* File: /media/ntfsdrive1/workspace/synchronizerchip/runset_pex/fullsystem_extracted.sp
* Created: Wed Dec  9 13:59:48 2015
* Program "Calibre xRC"
* Version "v2013.3_28.19"
* 
.include "/media/ntfsdrive1/workspace/synchronizerchip/runset_pex/fullsystem_extracted.sp.pex"
.subckt FULLSYSTEM 
* 
M0 45 N_12_M0_g N_32_M0_s N_32_X189/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=7e-14
+ AS=5.25e-14 PD=1.28e-06 PS=1.21e-06
M1 N_20_M1_d N_13_M1_g 45 N_32_X189/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=7e-14
+ AS=7e-14 PD=1.28e-06 PS=1.28e-06
M2 46 N_14_M2_g N_20_M1_d N_32_X189/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=7e-14
+ AS=7e-14 PD=1.28e-06 PS=1.28e-06
M3 N_32_M3_d N_21_M3_g 46 N_32_X189/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14
+ AS=7e-14 PD=1.21e-06 PS=1.28e-06
M4 47 N_28_M4_g N_31_M4_s N_32_X189/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=7e-14
+ AS=5.25e-14 PD=1.28e-06 PS=1.21e-06
M5 N_32_M5_d N_16_M5_g 47 N_32_X189/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=1.175e-13
+ AS=7e-14 PD=1.47e-06 PS=1.28e-06
M6 N_32_M6_d N_21_M6_g N_33_M6_s N_32_X188/M0_b NMOS_VTL L=5e-08 W=5e-07
+ AD=1.225e-13 AS=5.25e-14 PD=1.515e-06 PS=1.21e-06
M7 N_17_M7_d N_31_M7_g N_32_M5_d N_32_X189/M0_b NMOS_VTL L=5e-08 W=5e-07
+ AD=5.25e-14 AS=1.175e-13 PD=1.21e-06 PS=1.47e-06
M8 48 N_21_M8_g N_32_M6_d N_32_X188/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=7e-14
+ AS=1.225e-13 PD=1.28e-06 PS=1.515e-06
M9 N_16_M9_d N_19_M9_g 48 N_32_X188/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=7e-14
+ AS=7e-14 PD=1.28e-06 PS=1.28e-06
M10 49 N_36_M10_g N_16_M9_d N_32_X188/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=7e-14
+ AS=7e-14 PD=1.28e-06 PS=1.28e-06
M11 N_32_M11_d N_33_M11_g 49 N_32_X188/M0_b NMOS_VTL L=5e-08 W=5e-07
+ AD=2.025e-13 AS=7e-14 PD=1.81e-06 PS=1.28e-06
M12 N_34_M12_d N_19_M12_g N_32_M12_s N_32_X192/M0_b NMOS_VTL L=5e-08 W=2.5e-07
+ AD=3.5e-14 AS=2.625e-14 PD=7.8e-07 PS=7.1e-07
M13 N_32_M13_d N_20_M13_g N_34_M12_d N_32_X192/M0_b NMOS_VTL L=5e-08 W=2.5e-07
+ AD=7.875e-14 AS=3.5e-14 PD=1.49e-06 PS=7.8e-07
M14 N_36_M14_d N_19_M14_g N_32_M11_d N_32_X188/M0_b NMOS_VTL L=5e-08 W=5e-07
+ AD=5.25e-14 AS=2.025e-13 PD=1.21e-06 PS=1.81e-06
M15 N_37_M15_d N_34_M15_g N_32_M13_d N_32_X192/M0_b NMOS_VTL L=5e-08 W=5e-07
+ AD=5.25e-14 AS=7.875e-14 PD=1.21e-06 PS=1.49e-06
M16 N_38_M16_d N_21_M16_g N_32_M16_s N_32_X188/M0_b NMOS_VTL L=5e-08 W=2.5e-07
+ AD=3.5e-14 AS=2.625e-14 PD=7.8e-07 PS=7.1e-07
M17 N_32_M17_d N_16_M17_g N_38_M16_d N_32_X188/M0_b NMOS_VTL L=5e-08 W=2.5e-07
+ AD=2.625e-14 AS=3.5e-14 PD=7.1e-07 PS=7.8e-07
M18 N_20_M18_d N_12_M18_g N_30_M18_s N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.4e-13 AS=1.05e-13 PD=2.28e-06 PS=2.21e-06
M19 N_30_M19_d N_13_M19_g N_20_M18_d N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.4e-13 AS=1.4e-13 PD=2.28e-06 PS=2.28e-06
M20 N_22_M20_d N_14_M20_g N_30_M19_d N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.4e-13 AS=1.4e-13 PD=2.28e-06 PS=2.28e-06
M21 N_30_M21_d N_21_M21_g N_22_M20_d N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.05e-13 AS=1.4e-13 PD=2.21e-06 PS=2.28e-06
M22 N_31_M22_d N_28_M22_g N_22_M22_s N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07
+ AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.21e-06
M23 N_22_M23_d N_16_M23_g N_31_M22_d N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07
+ AD=1.575e-13 AS=7e-14 PD=2.49e-06 PS=1.28e-06
M24 N_22_M24_d N_21_M24_g N_33_M24_s N_22_X188/M1_b PMOS_VTL L=5e-08 W=1e-06
+ AD=3.05e-13 AS=1.05e-13 PD=2.61e-06 PS=2.21e-06
M25 N_17_M25_d N_31_M25_g N_22_M23_d N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.05e-13 AS=1.575e-13 PD=2.21e-06 PS=2.49e-06
M26 41 N_21_M26_g N_22_M24_d N_22_X188/M1_b PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13
+ AS=3.05e-13 PD=2.28e-06 PS=2.61e-06
M27 N_16_M27_d N_36_M27_g 41 N_22_X188/M1_b PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13
+ AS=1.4e-13 PD=2.28e-06 PS=2.28e-06
M28 42 N_19_M28_g N_16_M27_d N_22_X188/M1_b PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13
+ AS=1.4e-13 PD=2.28e-06 PS=2.28e-06
M29 43 N_19_M29_g N_34_M29_s N_22_X189/M1_b PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13
+ AS=1.05e-13 PD=2.28e-06 PS=2.21e-06
M30 N_22_M30_d N_33_M30_g 42 N_22_X188/M1_b PMOS_VTL L=5e-08 W=1e-06 AD=3.45e-13
+ AS=1.4e-13 PD=2.69e-06 PS=2.28e-06
M31 N_22_M31_d N_20_M31_g 43 N_22_X189/M1_b PMOS_VTL L=5e-08 W=1e-06 AD=2.45e-13
+ AS=1.4e-13 PD=2.49e-06 PS=2.28e-06
M32 N_36_M32_d N_19_M32_g N_22_M30_d N_22_X188/M1_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.05e-13 AS=3.45e-13 PD=2.21e-06 PS=2.69e-06
M33 N_37_M33_d N_34_M33_g N_22_M31_d N_22_X189/M1_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.05e-13 AS=2.45e-13 PD=2.21e-06 PS=2.49e-06
M34 44 N_21_M34_g N_22_M34_s N_22_X188/M1_b PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13
+ AS=1.05e-13 PD=2.28e-06 PS=2.21e-06
M35 N_38_M35_d N_16_M35_g 44 N_22_X188/M1_b PMOS_VTL L=5e-08 W=1e-06 AD=1.05e-13
+ AS=1.4e-13 PD=2.21e-06 PS=2.28e-06
mX188/M0 N_2_X188/M0_d N_23_X188/M0_g N_32_X188/M0_s N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX188/M1 N_2_X188/M1_d N_23_X188/M1_g N_22_X188/M1_s N_22_X188/M1_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX189/M0 N_24_X189/M0_d N_7_X189/M0_g N_32_X189/M0_s N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX189/M1 N_24_X189/M1_d N_7_X189/M1_g N_22_X189/M1_s N_22_X189/M1_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX190/M0 N_3_X190/M0_d N_25_X190/M0_g N_32_X190/M0_s N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX190/M1 N_3_X190/M1_d N_25_X190/M1_g N_22_X190/M1_s N_22_X188/M1_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX191/M0 N_25_X191/M0_d N_6_X191/M0_g N_32_X191/M0_s N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX191/M1 N_25_X191/M1_d N_6_X191/M1_g N_22_X191/M1_s N_22_X188/M1_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX192/M0 N_26_X192/M0_d N_9_X192/M0_g N_32_X192/M0_s N_32_X192/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX192/M1 N_26_X192/M1_d N_9_X192/M1_g N_22_X192/M1_s N_22_X192/M1_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX193/M0 N_14_X193/M0_d N_28_X193/M0_g N_32_X193/M0_s N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX193/M1 N_14_X193/M1_d N_28_X193/M1_g N_22_X193/M1_s N_22_X189/M1_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX194/X1/M0 N_23_X194/X1/M0_d N_15_X194/X1/M0_g N_32_X194/X1/M0_s N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX194/X1/M1 N_23_X194/X1/M1_d N_15_X194/X1/M1_g N_22_X194/X1/M1_s N_22_X188/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX195/X1/M0 N_5_X195/X1/M0_d N_24_X195/X1/M0_g N_32_X195/X1/M0_s N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX195/X1/M1 N_5_X195/X1/M1_d N_24_X195/X1/M1_g N_22_X195/X1/M1_s N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX196/X1/M0 N_8_X196/X1/M0_d N_26_X196/X1/M0_g N_32_X196/X1/M0_s N_32_X192/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX196/X1/M1 N_8_X196/X1/M1_d N_26_X196/X1/M1_g N_22_X196/X1/M1_s N_22_X192/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX197/X1/M0 N_10_X197/X1/M0_d N_27_X197/X1/M0_g N_32_X197/X1/M0_s N_32_X192/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX197/X1/M1 N_10_X197/X1/M1_d N_27_X197/X1/M1_g N_22_X197/X1/M1_s N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX198/X1/M0 N_13_X198/X1/M0_d N_21_X198/X1/M0_g N_32_X198/X1/M0_s N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX198/X1/M1 N_13_X198/X1/M1_d N_21_X198/X1/M1_g N_22_X198/X1/M1_s
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06
+ PS=1.21e-06
mX199/X1/M0 N_27_X199/X1/M0_d N_18_X199/X1/M0_g N_32_X199/X1/M0_s N_32_X192/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX199/X1/M1 N_27_X199/X1/M1_d N_18_X199/X1/M1_g N_22_X199/X1/M1_s N_22_X192/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX200/X1/M0 N_29_X200/X1/M0_d N_39_X200/X1/M0_g N_32_X200/X1/M0_s N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX200/X1/M1 N_29_X200/X1/M1_d N_39_X200/X1/M1_g N_22_X200/X1/M1_s N_22_X188/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX201/X1/M0 N_35_X201/X1/M0_d N_40_X201/X1/M0_g N_32_X201/X1/M0_s N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX201/X1/M1 N_35_X201/X1/M1_d N_40_X201/X1/M1_g N_22_X201/X1/M1_s
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06
+ PS=1.21e-06
mX202/X1/M0 N_11_X202/X1/M0_d N_37_X202/X1/M0_g N_32_X202/X1/M0_s N_32_X192/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX202/X1/M1 N_11_X202/X1/M1_d N_37_X202/X1/M1_g N_22_X202/X1/M1_s N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX203/M0 N_32_X203/M0_d N_1_X203/M0_g N_X203/10_X203/M0_s N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX203/M1 N_X203/11_X203/M1_d N_2_X203/M1_g N_32_X203/M0_d N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX203/M2 N_X203/9_X203/M2_d N_X203/10_X203/M2_g N_32_X203/M2_s N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX203/M3 N_X203/13_X203/M3_d N_X203/10_X203/M3_g N_X203/11_X203/M1_d
+ N_32_X188/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06
+ PS=9.2e-07
mX203/M4 N_X203/12_X203/M4_d N_X203/9_X203/M4_g N_X203/13_X203/M3_d
+ N_32_X188/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06
+ PS=1.2e-06
mX203/M5 X203/18 N_29_X203/M5_g N_X203/12_X203/M4_d N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX203/M6 N_32_X203/M6_d N_X203/14_X203/M6_g X203/18 N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX203/M7 X203/19 N_X203/13_X203/M7_g N_32_X203/M6_d N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX203/M8 N_X203/14_X203/M8_d N_22_X203/M8_g X203/19 N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX203/M9 N_X203/16_X203/M9_d N_X203/9_X203/M9_g N_X203/14_X203/M8_d
+ N_32_X188/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06
+ PS=1.38e-06
mX203/M10 N_X203/15_X203/M10_d N_X203/10_X203/M10_g N_X203/16_X203/M9_d
+ N_32_X188/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06
+ PS=1.04e-06
mX203/M11 X203/20 N_22_X203/M11_g N_X203/15_X203/M10_d N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX203/M12 N_32_X203/M12_d N_X203/17_X203/M12_g X203/20 N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX203/M13 X203/21 N_29_X203/M13_g N_32_X203/M12_d N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX203/M14 N_X203/17_X203/M14_d N_X203/16_X203/M14_g X203/21 N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX203/M15 N_6_X203/M15_d N_X203/17_X203/M15_g N_32_X203/M15_s N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX203/M16 N_22_X203/M16_d N_1_X203/M16_g N_X203/10_X203/M16_s N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX203/M17 N_X203/11_X203/M17_d N_2_X203/M17_g N_22_X203/M16_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX203/M18 N_X203/13_X203/M18_d N_X203/9_X203/M18_g N_X203/11_X203/M17_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14
+ PD=1.09e-06 PS=1.28e-06
mX203/M19 N_X203/12_X203/M19_d N_X203/10_X203/M19_g N_X203/13_X203/M18_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14
+ PD=1.38e-06 PS=1.09e-06
mX203/M20 N_22_X203/M20_d N_X203/10_X203/M20_g N_X203/9_X203/M20_s
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06
+ PS=1.21e-06
mX203/M21 N_22_X203/M21_d N_29_X203/M21_g N_X203/12_X203/M19_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX203/M22 N_X203/12_X203/M22_d N_X203/14_X203/M22_g N_22_X203/M21_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13
+ PD=1.21e-06 PS=2.33e-06
mX203/M23 N_X203/14_X203/M23_d N_22_X203/M23_g N_22_X203/M23_s N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX203/M24 N_X203/16_X203/M24_d N_X203/10_X203/M24_g N_X203/14_X203/M23_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13
+ PD=7.8e-07 PS=3.12e-06
mX203/M25 N_22_X203/M25_d N_X203/13_X203/M25_g N_X203/14_X203/M23_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX203/M26 N_X203/15_X203/M26_d N_X203/9_X203/M26_g N_X203/16_X203/M24_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14
+ PD=3.3e-06 PS=7.8e-07
mX203/M27 N_X203/15_X203/M26_d N_X203/17_X203/M27_g N_22_X203/M25_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX203/M28 N_22_X203/M28_d N_22_X203/M28_g N_X203/15_X203/M26_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX203/M29 N_X203/17_X203/M29_d N_29_X203/M29_g N_22_X203/M28_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX203/M30 N_22_X203/M30_d N_X203/16_X203/M30_g N_X203/17_X203/M29_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06
+ PS=1.28e-06
mX203/M31 N_6_X203/M31_d N_X203/17_X203/M31_g N_22_X203/M30_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
mX204/M0 N_32_X204/M0_d N_1_X204/M0_g N_X204/10_X204/M0_s N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX204/M1 N_X204/11_X204/M1_d N_3_X204/M1_g N_32_X204/M0_d N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX204/M2 N_X204/9_X204/M2_d N_X204/10_X204/M2_g N_32_X204/M2_s N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX204/M3 N_X204/13_X204/M3_d N_X204/10_X204/M3_g N_X204/11_X204/M1_d
+ N_32_X189/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06
+ PS=9.2e-07
mX204/M4 N_X204/12_X204/M4_d N_X204/9_X204/M4_g N_X204/13_X204/M3_d
+ N_32_X189/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06
+ PS=1.2e-06
mX204/M5 X204/18 N_29_X204/M5_g N_X204/12_X204/M4_d N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX204/M6 N_32_X204/M6_d N_X204/14_X204/M6_g X204/18 N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX204/M7 X204/19 N_X204/13_X204/M7_g N_32_X204/M6_d N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX204/M8 N_X204/14_X204/M8_d N_22_X204/M8_g X204/19 N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX204/M9 N_X204/16_X204/M9_d N_X204/9_X204/M9_g N_X204/14_X204/M8_d
+ N_32_X189/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06
+ PS=1.38e-06
mX204/M10 N_X204/15_X204/M10_d N_X204/10_X204/M10_g N_X204/16_X204/M9_d
+ N_32_X189/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06
+ PS=1.04e-06
mX204/M11 X204/20 N_22_X204/M11_g N_X204/15_X204/M10_d N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX204/M12 N_32_X204/M12_d N_X204/17_X204/M12_g X204/20 N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX204/M13 X204/21 N_29_X204/M13_g N_32_X204/M12_d N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX204/M14 N_X204/17_X204/M14_d N_X204/16_X204/M14_g X204/21 N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX204/M15 N_7_X204/M15_d N_X204/17_X204/M15_g N_32_X204/M15_s N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX204/M16 N_22_X204/M16_d N_1_X204/M16_g N_X204/10_X204/M16_s N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX204/M17 N_X204/11_X204/M17_d N_3_X204/M17_g N_22_X204/M16_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX204/M18 N_X204/13_X204/M18_d N_X204/9_X204/M18_g N_X204/11_X204/M17_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14
+ PD=1.09e-06 PS=1.28e-06
mX204/M19 N_X204/12_X204/M19_d N_X204/10_X204/M19_g N_X204/13_X204/M18_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14
+ PD=1.38e-06 PS=1.09e-06
mX204/M20 N_22_X204/M20_d N_X204/10_X204/M20_g N_X204/9_X204/M20_s
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06
+ PS=1.21e-06
mX204/M21 N_22_X204/M21_d N_29_X204/M21_g N_X204/12_X204/M19_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX204/M22 N_X204/12_X204/M22_d N_X204/14_X204/M22_g N_22_X204/M21_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13
+ PD=1.21e-06 PS=2.33e-06
mX204/M23 N_X204/14_X204/M23_d N_22_X204/M23_g N_22_X204/M23_s N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX204/M24 N_X204/16_X204/M24_d N_X204/10_X204/M24_g N_X204/14_X204/M23_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13
+ PD=7.8e-07 PS=3.12e-06
mX204/M25 N_22_X204/M25_d N_X204/13_X204/M25_g N_X204/14_X204/M23_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX204/M26 N_X204/15_X204/M26_d N_X204/9_X204/M26_g N_X204/16_X204/M24_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14
+ PD=3.3e-06 PS=7.8e-07
mX204/M27 N_X204/15_X204/M26_d N_X204/17_X204/M27_g N_22_X204/M25_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX204/M28 N_22_X204/M28_d N_22_X204/M28_g N_X204/15_X204/M26_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX204/M29 N_X204/17_X204/M29_d N_29_X204/M29_g N_22_X204/M28_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX204/M30 N_22_X204/M30_d N_X204/16_X204/M30_g N_X204/17_X204/M29_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06
+ PS=1.28e-06
mX204/M31 N_7_X204/M31_d N_X204/17_X204/M31_g N_22_X204/M30_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
mX205/M0 N_32_X205/M0_d N_4_X205/M0_g N_X205/10_X205/M0_s N_32_X192/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX205/M1 N_X205/11_X205/M1_d N_5_X205/M1_g N_32_X205/M0_d N_32_X192/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX205/M2 N_X205/9_X205/M2_d N_X205/10_X205/M2_g N_32_X205/M2_s N_32_X192/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX205/M3 N_X205/13_X205/M3_d N_X205/10_X205/M3_g N_X205/11_X205/M1_d
+ N_32_X192/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06
+ PS=9.2e-07
mX205/M4 N_X205/12_X205/M4_d N_X205/9_X205/M4_g N_X205/13_X205/M3_d
+ N_32_X192/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06
+ PS=1.2e-06
mX205/M5 X205/18 N_35_X205/M5_g N_X205/12_X205/M4_d N_32_X192/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX205/M6 N_32_X205/M6_d N_X205/14_X205/M6_g X205/18 N_32_X192/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX205/M7 X205/19 N_X205/13_X205/M7_g N_32_X205/M6_d N_32_X192/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX205/M8 N_X205/14_X205/M8_d N_22_X205/M8_g X205/19 N_32_X192/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX205/M9 N_X205/16_X205/M9_d N_X205/9_X205/M9_g N_X205/14_X205/M8_d
+ N_32_X192/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06
+ PS=1.38e-06
mX205/M10 N_X205/15_X205/M10_d N_X205/10_X205/M10_g N_X205/16_X205/M9_d
+ N_32_X192/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06
+ PS=1.04e-06
mX205/M11 X205/20 N_22_X205/M11_g N_X205/15_X205/M10_d N_32_X192/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX205/M12 N_32_X205/M12_d N_X205/17_X205/M12_g X205/20 N_32_X192/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX205/M13 X205/21 N_35_X205/M13_g N_32_X205/M12_d N_32_X192/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX205/M14 N_X205/17_X205/M14_d N_X205/16_X205/M14_g X205/21 N_32_X192/M0_b
+ NMOS_VTL L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX205/M15 N_9_X205/M15_d N_X205/17_X205/M15_g N_32_X205/M15_s N_32_X192/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX205/M16 N_22_X205/M16_d N_4_X205/M16_g N_X205/10_X205/M16_s N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX205/M17 N_X205/11_X205/M17_d N_5_X205/M17_g N_22_X205/M16_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX205/M18 N_X205/13_X205/M18_d N_X205/9_X205/M18_g N_X205/11_X205/M17_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14 PD=1.09e-06
+ PS=1.28e-06
mX205/M19 N_X205/12_X205/M19_d N_X205/10_X205/M19_g N_X205/13_X205/M18_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14 PD=1.38e-06
+ PS=1.09e-06
mX205/M20 N_22_X205/M20_d N_X205/10_X205/M20_g N_X205/9_X205/M20_s
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06
+ PS=1.21e-06
mX205/M21 N_22_X205/M21_d N_35_X205/M21_g N_X205/12_X205/M19_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX205/M22 N_X205/12_X205/M22_d N_X205/14_X205/M22_g N_22_X205/M21_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13 PD=1.21e-06
+ PS=2.33e-06
mX205/M23 N_X205/14_X205/M23_d N_22_X205/M23_g N_22_X205/M23_s N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX205/M24 N_X205/16_X205/M24_d N_X205/10_X205/M24_g N_X205/14_X205/M23_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13 PD=7.8e-07
+ PS=3.12e-06
mX205/M25 N_22_X205/M25_d N_X205/13_X205/M25_g N_X205/14_X205/M23_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX205/M26 N_X205/15_X205/M26_d N_X205/9_X205/M26_g N_X205/16_X205/M24_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14 PD=3.3e-06
+ PS=7.8e-07
mX205/M27 N_X205/15_X205/M26_d N_X205/17_X205/M27_g N_22_X205/M25_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX205/M28 N_22_X205/M28_d N_22_X205/M28_g N_X205/15_X205/M26_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX205/M29 N_X205/17_X205/M29_d N_35_X205/M29_g N_22_X205/M28_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX205/M30 N_22_X205/M30_d N_X205/16_X205/M30_g N_X205/17_X205/M29_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06
+ PS=1.28e-06
mX205/M31 N_9_X205/M31_d N_X205/17_X205/M31_g N_22_X205/M30_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
mX206/M0 N_32_X206/M0_d N_4_X206/M0_g N_X206/10_X206/M0_s N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX206/M1 N_X206/11_X206/M1_d N_8_X206/M1_g N_32_X206/M0_d N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX206/M2 N_X206/9_X206/M2_d N_X206/10_X206/M2_g N_32_X206/M2_s N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX206/M3 N_X206/13_X206/M3_d N_X206/10_X206/M3_g N_X206/11_X206/M1_d
+ N_32_X189/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06
+ PS=9.2e-07
mX206/M4 N_X206/12_X206/M4_d N_X206/9_X206/M4_g N_X206/13_X206/M3_d
+ N_32_X189/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06
+ PS=1.2e-06
mX206/M5 X206/18 N_35_X206/M5_g N_X206/12_X206/M4_d N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX206/M6 N_32_X206/M6_d N_X206/14_X206/M6_g X206/18 N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX206/M7 X206/19 N_X206/13_X206/M7_g N_32_X206/M6_d N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX206/M8 N_X206/14_X206/M8_d N_22_X206/M8_g X206/19 N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX206/M9 N_X206/16_X206/M9_d N_X206/9_X206/M9_g N_X206/14_X206/M8_d
+ N_32_X189/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06
+ PS=1.38e-06
mX206/M10 N_X206/15_X206/M10_d N_X206/10_X206/M10_g N_X206/16_X206/M9_d
+ N_32_X189/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06
+ PS=1.04e-06
mX206/M11 X206/20 N_22_X206/M11_g N_X206/15_X206/M10_d N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX206/M12 N_32_X206/M12_d N_X206/17_X206/M12_g X206/20 N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX206/M13 X206/21 N_35_X206/M13_g N_32_X206/M12_d N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX206/M14 N_X206/17_X206/M14_d N_X206/16_X206/M14_g X206/21 N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX206/M15 N_28_X206/M15_d N_X206/17_X206/M15_g N_32_X206/M15_s N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX206/M16 N_22_X206/M16_d N_4_X206/M16_g N_X206/10_X206/M16_s N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX206/M17 N_X206/11_X206/M17_d N_8_X206/M17_g N_22_X206/M16_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX206/M18 N_X206/13_X206/M18_d N_X206/9_X206/M18_g N_X206/11_X206/M17_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14 PD=1.09e-06
+ PS=1.28e-06
mX206/M19 N_X206/12_X206/M19_d N_X206/10_X206/M19_g N_X206/13_X206/M18_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14 PD=1.38e-06
+ PS=1.09e-06
mX206/M20 N_22_X206/M20_d N_X206/10_X206/M20_g N_X206/9_X206/M20_s
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06
+ PS=1.21e-06
mX206/M21 N_22_X206/M21_d N_35_X206/M21_g N_X206/12_X206/M19_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX206/M22 N_X206/12_X206/M22_d N_X206/14_X206/M22_g N_22_X206/M21_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13 PD=1.21e-06
+ PS=2.33e-06
mX206/M23 N_X206/14_X206/M23_d N_22_X206/M23_g N_22_X206/M23_s N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX206/M24 N_X206/16_X206/M24_d N_X206/10_X206/M24_g N_X206/14_X206/M23_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13 PD=7.8e-07
+ PS=3.12e-06
mX206/M25 N_22_X206/M25_d N_X206/13_X206/M25_g N_X206/14_X206/M23_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX206/M26 N_X206/15_X206/M26_d N_X206/9_X206/M26_g N_X206/16_X206/M24_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14 PD=3.3e-06
+ PS=7.8e-07
mX206/M27 N_X206/15_X206/M26_d N_X206/17_X206/M27_g N_22_X206/M25_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX206/M28 N_22_X206/M28_d N_22_X206/M28_g N_X206/15_X206/M26_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX206/M29 N_X206/17_X206/M29_d N_35_X206/M29_g N_22_X206/M28_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX206/M30 N_22_X206/M30_d N_X206/16_X206/M30_g N_X206/17_X206/M29_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06
+ PS=1.28e-06
mX206/M31 N_28_X206/M31_d N_X206/17_X206/M31_g N_22_X206/M30_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
mX207/M0 N_32_X207/M0_d N_1_X207/M0_g N_X207/10_X207/M0_s N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX207/M1 N_X207/11_X207/M1_d N_10_X207/M1_g N_32_X207/M0_d N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX207/M2 N_X207/9_X207/M2_d N_X207/10_X207/M2_g N_32_X207/M2_s N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX207/M3 N_X207/13_X207/M3_d N_X207/10_X207/M3_g N_X207/11_X207/M1_d
+ N_32_X188/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06
+ PS=9.2e-07
mX207/M4 N_X207/12_X207/M4_d N_X207/9_X207/M4_g N_X207/13_X207/M3_d
+ N_32_X188/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06
+ PS=1.2e-06
mX207/M5 X207/18 N_29_X207/M5_g N_X207/12_X207/M4_d N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX207/M6 N_32_X207/M6_d N_X207/14_X207/M6_g X207/18 N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX207/M7 X207/19 N_X207/13_X207/M7_g N_32_X207/M6_d N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX207/M8 N_X207/14_X207/M8_d N_22_X207/M8_g X207/19 N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX207/M9 N_X207/16_X207/M9_d N_X207/9_X207/M9_g N_X207/14_X207/M8_d
+ N_32_X188/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06
+ PS=1.38e-06
mX207/M10 N_X207/15_X207/M10_d N_X207/10_X207/M10_g N_X207/16_X207/M9_d
+ N_32_X188/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06
+ PS=1.04e-06
mX207/M11 X207/20 N_22_X207/M11_g N_X207/15_X207/M10_d N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX207/M12 N_32_X207/M12_d N_X207/17_X207/M12_g X207/20 N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX207/M13 X207/21 N_29_X207/M13_g N_32_X207/M12_d N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX207/M14 N_X207/17_X207/M14_d N_X207/16_X207/M14_g X207/21 N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX207/M15 N_15_X207/M15_d N_X207/17_X207/M15_g N_32_X207/M15_s N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX207/M16 N_22_X207/M16_d N_1_X207/M16_g N_X207/10_X207/M16_s N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX207/M17 N_X207/11_X207/M17_d N_10_X207/M17_g N_22_X207/M16_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX207/M18 N_X207/13_X207/M18_d N_X207/9_X207/M18_g N_X207/11_X207/M17_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14
+ PD=1.09e-06 PS=1.28e-06
mX207/M19 N_X207/12_X207/M19_d N_X207/10_X207/M19_g N_X207/13_X207/M18_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14
+ PD=1.38e-06 PS=1.09e-06
mX207/M20 N_22_X207/M20_d N_X207/10_X207/M20_g N_X207/9_X207/M20_s
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06
+ PS=1.21e-06
mX207/M21 N_22_X207/M21_d N_29_X207/M21_g N_X207/12_X207/M19_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX207/M22 N_X207/12_X207/M22_d N_X207/14_X207/M22_g N_22_X207/M21_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13
+ PD=1.21e-06 PS=2.33e-06
mX207/M23 N_X207/14_X207/M23_d N_22_X207/M23_g N_22_X207/M23_s N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX207/M24 N_X207/16_X207/M24_d N_X207/10_X207/M24_g N_X207/14_X207/M23_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13
+ PD=7.8e-07 PS=3.12e-06
mX207/M25 N_22_X207/M25_d N_X207/13_X207/M25_g N_X207/14_X207/M23_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX207/M26 N_X207/15_X207/M26_d N_X207/9_X207/M26_g N_X207/16_X207/M24_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14
+ PD=3.3e-06 PS=7.8e-07
mX207/M27 N_X207/15_X207/M26_d N_X207/17_X207/M27_g N_22_X207/M25_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX207/M28 N_22_X207/M28_d N_22_X207/M28_g N_X207/15_X207/M26_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX207/M29 N_X207/17_X207/M29_d N_29_X207/M29_g N_22_X207/M28_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX207/M30 N_22_X207/M30_d N_X207/16_X207/M30_g N_X207/17_X207/M29_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06
+ PS=1.28e-06
mX207/M31 N_15_X207/M31_d N_X207/17_X207/M31_g N_22_X207/M30_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
mX208/M0 N_32_X208/M0_d N_4_X208/M0_g N_X208/10_X208/M0_s N_32_X192/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX208/M1 N_X208/11_X208/M1_d N_11_X208/M1_g N_32_X208/M0_d N_32_X192/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX208/M2 N_X208/9_X208/M2_d N_X208/10_X208/M2_g N_32_X208/M2_s N_32_X192/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX208/M3 N_X208/13_X208/M3_d N_X208/10_X208/M3_g N_X208/11_X208/M1_d
+ N_32_X192/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06
+ PS=9.2e-07
mX208/M4 N_X208/12_X208/M4_d N_X208/9_X208/M4_g N_X208/13_X208/M3_d
+ N_32_X192/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06
+ PS=1.2e-06
mX208/M5 X208/18 N_35_X208/M5_g N_X208/12_X208/M4_d N_32_X192/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX208/M6 N_32_X208/M6_d N_X208/14_X208/M6_g X208/18 N_32_X192/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX208/M7 X208/19 N_X208/13_X208/M7_g N_32_X208/M6_d N_32_X192/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX208/M8 N_X208/14_X208/M8_d N_22_X208/M8_g X208/19 N_32_X192/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX208/M9 N_X208/16_X208/M9_d N_X208/9_X208/M9_g N_X208/14_X208/M8_d
+ N_32_X192/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06
+ PS=1.38e-06
mX208/M10 N_X208/15_X208/M10_d N_X208/10_X208/M10_g N_X208/16_X208/M9_d
+ N_32_X192/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06
+ PS=1.04e-06
mX208/M11 X208/20 N_22_X208/M11_g N_X208/15_X208/M10_d N_32_X192/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX208/M12 N_32_X208/M12_d N_X208/17_X208/M12_g X208/20 N_32_X192/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX208/M13 X208/21 N_35_X208/M13_g N_32_X208/M12_d N_32_X192/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX208/M14 N_X208/17_X208/M14_d N_X208/16_X208/M14_g X208/21 N_32_X192/M0_b
+ NMOS_VTL L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX208/M15 N_18_X208/M15_d N_X208/17_X208/M15_g N_32_X208/M15_s N_32_X192/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX208/M16 N_22_X208/M16_d N_4_X208/M16_g N_X208/10_X208/M16_s N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX208/M17 N_X208/11_X208/M17_d N_11_X208/M17_g N_22_X208/M16_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX208/M18 N_X208/13_X208/M18_d N_X208/9_X208/M18_g N_X208/11_X208/M17_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14 PD=1.09e-06
+ PS=1.28e-06
mX208/M19 N_X208/12_X208/M19_d N_X208/10_X208/M19_g N_X208/13_X208/M18_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14 PD=1.38e-06
+ PS=1.09e-06
mX208/M20 N_22_X208/M20_d N_X208/10_X208/M20_g N_X208/9_X208/M20_s
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06
+ PS=1.21e-06
mX208/M21 N_22_X208/M21_d N_35_X208/M21_g N_X208/12_X208/M19_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX208/M22 N_X208/12_X208/M22_d N_X208/14_X208/M22_g N_22_X208/M21_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13 PD=1.21e-06
+ PS=2.33e-06
mX208/M23 N_X208/14_X208/M23_d N_22_X208/M23_g N_22_X208/M23_s N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX208/M24 N_X208/16_X208/M24_d N_X208/10_X208/M24_g N_X208/14_X208/M23_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13 PD=7.8e-07
+ PS=3.12e-06
mX208/M25 N_22_X208/M25_d N_X208/13_X208/M25_g N_X208/14_X208/M23_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX208/M26 N_X208/15_X208/M26_d N_X208/9_X208/M26_g N_X208/16_X208/M24_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14 PD=3.3e-06
+ PS=7.8e-07
mX208/M27 N_X208/15_X208/M26_d N_X208/17_X208/M27_g N_22_X208/M25_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX208/M28 N_22_X208/M28_d N_22_X208/M28_g N_X208/15_X208/M26_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX208/M29 N_X208/17_X208/M29_d N_35_X208/M29_g N_22_X208/M28_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX208/M30 N_22_X208/M30_d N_X208/16_X208/M30_g N_X208/17_X208/M29_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06
+ PS=1.28e-06
mX208/M31 N_18_X208/M31_d N_X208/17_X208/M31_g N_22_X208/M30_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
mX209/M0 N_32_X209/M0_d N_4_X209/M0_g N_X209/10_X209/M0_s N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX209/M1 N_X209/11_X209/M1_d N_11_X209/M1_g N_32_X209/M0_d N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX209/M2 N_X209/9_X209/M2_d N_X209/10_X209/M2_g N_32_X209/M2_s N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX209/M3 N_X209/13_X209/M3_d N_X209/10_X209/M3_g N_X209/11_X209/M1_d
+ N_32_X189/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06
+ PS=9.2e-07
mX209/M4 N_X209/12_X209/M4_d N_X209/9_X209/M4_g N_X209/13_X209/M3_d
+ N_32_X189/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06
+ PS=1.2e-06
mX209/M5 X209/18 N_35_X209/M5_g N_X209/12_X209/M4_d N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX209/M6 N_32_X209/M6_d N_X209/14_X209/M6_g X209/18 N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX209/M7 X209/19 N_X209/13_X209/M7_g N_32_X209/M6_d N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX209/M8 N_X209/14_X209/M8_d N_22_X209/M8_g X209/19 N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX209/M9 N_X209/16_X209/M9_d N_X209/9_X209/M9_g N_X209/14_X209/M8_d
+ N_32_X189/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06
+ PS=1.38e-06
mX209/M10 N_X209/15_X209/M10_d N_X209/10_X209/M10_g N_X209/16_X209/M9_d
+ N_32_X189/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06
+ PS=1.04e-06
mX209/M11 X209/20 N_22_X209/M11_g N_X209/15_X209/M10_d N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX209/M12 N_32_X209/M12_d N_X209/17_X209/M12_g X209/20 N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX209/M13 X209/21 N_35_X209/M13_g N_32_X209/M12_d N_32_X189/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX209/M14 N_X209/17_X209/M14_d N_X209/16_X209/M14_g X209/21 N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX209/M15 N_21_X209/M15_d N_X209/17_X209/M15_g N_32_X209/M15_s N_32_X189/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX209/M16 N_22_X209/M16_d N_4_X209/M16_g N_X209/10_X209/M16_s N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX209/M17 N_X209/11_X209/M17_d N_11_X209/M17_g N_22_X209/M16_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX209/M18 N_X209/13_X209/M18_d N_X209/9_X209/M18_g N_X209/11_X209/M17_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14 PD=1.09e-06
+ PS=1.28e-06
mX209/M19 N_X209/12_X209/M19_d N_X209/10_X209/M19_g N_X209/13_X209/M18_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14 PD=1.38e-06
+ PS=1.09e-06
mX209/M20 N_22_X209/M20_d N_X209/10_X209/M20_g N_X209/9_X209/M20_s
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06
+ PS=1.21e-06
mX209/M21 N_22_X209/M21_d N_35_X209/M21_g N_X209/12_X209/M19_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX209/M22 N_X209/12_X209/M22_d N_X209/14_X209/M22_g N_22_X209/M21_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13 PD=1.21e-06
+ PS=2.33e-06
mX209/M23 N_X209/14_X209/M23_d N_22_X209/M23_g N_22_X209/M23_s N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX209/M24 N_X209/16_X209/M24_d N_X209/10_X209/M24_g N_X209/14_X209/M23_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13 PD=7.8e-07
+ PS=3.12e-06
mX209/M25 N_22_X209/M25_d N_X209/13_X209/M25_g N_X209/14_X209/M23_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX209/M26 N_X209/15_X209/M26_d N_X209/9_X209/M26_g N_X209/16_X209/M24_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14 PD=3.3e-06
+ PS=7.8e-07
mX209/M27 N_X209/15_X209/M26_d N_X209/17_X209/M27_g N_22_X209/M25_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX209/M28 N_22_X209/M28_d N_22_X209/M28_g N_X209/15_X209/M26_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX209/M29 N_X209/17_X209/M29_d N_35_X209/M29_g N_22_X209/M28_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX209/M30 N_22_X209/M30_d N_X209/16_X209/M30_g N_X209/17_X209/M29_d
+ N_22_X189/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06
+ PS=1.28e-06
mX209/M31 N_21_X209/M31_d N_X209/17_X209/M31_g N_22_X209/M30_d N_22_X189/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
mX210/M0 N_32_X210/M0_d N_4_X210/M0_g N_X210/10_X210/M0_s N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX210/M1 N_X210/11_X210/M1_d N_17_X210/M1_g N_32_X210/M0_d N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX210/M2 N_X210/9_X210/M2_d N_X210/10_X210/M2_g N_32_X210/M2_s N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX210/M3 N_X210/13_X210/M3_d N_X210/10_X210/M3_g N_X210/11_X210/M1_d
+ N_32_X188/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06
+ PS=9.2e-07
mX210/M4 N_X210/12_X210/M4_d N_X210/9_X210/M4_g N_X210/13_X210/M3_d
+ N_32_X188/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06
+ PS=1.2e-06
mX210/M5 X210/18 N_35_X210/M5_g N_X210/12_X210/M4_d N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX210/M6 N_32_X210/M6_d N_X210/14_X210/M6_g X210/18 N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX210/M7 X210/19 N_X210/13_X210/M7_g N_32_X210/M6_d N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX210/M8 N_X210/14_X210/M8_d N_22_X210/M8_g X210/19 N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX210/M9 N_X210/16_X210/M9_d N_X210/9_X210/M9_g N_X210/14_X210/M8_d
+ N_32_X188/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06
+ PS=1.38e-06
mX210/M10 N_X210/15_X210/M10_d N_X210/10_X210/M10_g N_X210/16_X210/M9_d
+ N_32_X188/M0_b NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06
+ PS=1.04e-06
mX210/M11 X210/20 N_22_X210/M11_g N_X210/15_X210/M10_d N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX210/M12 N_32_X210/M12_d N_X210/17_X210/M12_g X210/20 N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX210/M13 X210/21 N_35_X210/M13_g N_32_X210/M12_d N_32_X188/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX210/M14 N_X210/17_X210/M14_d N_X210/16_X210/M14_g X210/21 N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX210/M15 N_19_X210/M15_d N_X210/17_X210/M15_g N_32_X210/M15_s N_32_X188/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX210/M16 N_22_X210/M16_d N_4_X210/M16_g N_X210/10_X210/M16_s N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX210/M17 N_X210/11_X210/M17_d N_17_X210/M17_g N_22_X210/M16_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX210/M18 N_X210/13_X210/M18_d N_X210/9_X210/M18_g N_X210/11_X210/M17_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14
+ PD=1.09e-06 PS=1.28e-06
mX210/M19 N_X210/12_X210/M19_d N_X210/10_X210/M19_g N_X210/13_X210/M18_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14
+ PD=1.38e-06 PS=1.09e-06
mX210/M20 N_22_X210/M20_d N_X210/10_X210/M20_g N_X210/9_X210/M20_s
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06
+ PS=1.21e-06
mX210/M21 N_22_X210/M21_d N_35_X210/M21_g N_X210/12_X210/M19_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX210/M22 N_X210/12_X210/M22_d N_X210/14_X210/M22_g N_22_X210/M21_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13
+ PD=1.21e-06 PS=2.33e-06
mX210/M23 N_X210/14_X210/M23_d N_22_X210/M23_g N_22_X210/M23_s N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX210/M24 N_X210/16_X210/M24_d N_X210/10_X210/M24_g N_X210/14_X210/M23_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13
+ PD=7.8e-07 PS=3.12e-06
mX210/M25 N_22_X210/M25_d N_X210/13_X210/M25_g N_X210/14_X210/M23_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX210/M26 N_X210/15_X210/M26_d N_X210/9_X210/M26_g N_X210/16_X210/M24_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14
+ PD=3.3e-06 PS=7.8e-07
mX210/M27 N_X210/15_X210/M26_d N_X210/17_X210/M27_g N_22_X210/M25_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX210/M28 N_22_X210/M28_d N_22_X210/M28_g N_X210/15_X210/M26_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX210/M29 N_X210/17_X210/M29_d N_35_X210/M29_g N_22_X210/M28_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX210/M30 N_22_X210/M30_d N_X210/16_X210/M30_g N_X210/17_X210/M29_d
+ N_22_X198/X1/M1_b PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06
+ PS=1.28e-06
mX210/M31 N_19_X210/M31_d N_X210/17_X210/M31_g N_22_X210/M30_d N_22_X198/X1/M1_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
*
.include "/media/ntfsdrive1/workspace/synchronizerchip/runset_pex/fullsystem_extracted.sp.FULLSYSTEM.pxi"
*
.ends
*
*
