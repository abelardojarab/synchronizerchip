* SPICE NETLIST
***************************************

.SUBCKT M6_M5_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M5_M4_3
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M4_M3_2
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M6_M5_4
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M3_M2_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M2_M1_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=5 FDC=0
.ENDS
***************************************
.SUBCKT M2_M1_via
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M3_M2_via
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILL
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT INVX1 A gnd vdd Y
** N=4 EP=4 IP=0 FDC=2
* PORT A A 415 1110 metal1
* PORT gnd gnd 390 490 metal1
* PORT vdd vdd 390 3670 metal1
* PORT Y Y 760 2030 metal1
M0 Y A gnd gnd NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07 $X=525 $Y=355 $D=1
M1 Y A vdd vdd PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06 $X=525 $Y=2580 $D=0
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4
** N=4 EP=4 IP=6 FDC=2
X1 3 1 2 4 INVX1 $T=760 0 0 0 $X=560 $Y=-200
.ENDS
***************************************
.SUBCKT DFFSR CLK D S R vdd gnd Q 8
** N=21 EP=8 IP=0 FDC=32
* PORT CLK CLK 760 2190 metal1
* PORT D D 1140 1800 metal1
* PORT S S 5335 1970 metal1
* PORT R R 4815 3835 metal1
* PORT vdd vdd 4140 4420 metal1
* PORT gnd gnd 3480 575 metal1
* PORT Q Q 8030 1890 metal1
M0 gnd CLK 10 gnd NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07 $X=645 $Y=1310 $D=1
M1 11 D gnd gnd NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07 $X=1165 $Y=1310 $D=1
M2 9 10 gnd gnd NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07 $X=1685 $Y=530 $D=1
M3 13 10 11 gnd NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06 PS=9.2e-07 $X=1685 $Y=1310 $D=1
M4 12 9 13 gnd NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06 PS=1.2e-06 $X=2485 $Y=1310 $D=1
M5 18 R 12 gnd NMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06 $X=2865 $Y=810 $D=1
M6 gnd 14 18 gnd NMOS_VTL L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06 $X=3245 $Y=810 $D=1
M7 19 13 gnd gnd NMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06 $X=4065 $Y=810 $D=1
M8 14 S 19 gnd NMOS_VTL L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06 $X=4445 $Y=810 $D=1
M9 16 9 14 gnd NMOS_VTL L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06 PS=1.38e-06 $X=4925 $Y=1100 $D=1
M10 15 10 16 gnd NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06 PS=1.04e-06 $X=5565 $Y=1100 $D=1
M11 20 S 15 gnd NMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06 $X=5945 $Y=600 $D=1
M12 gnd 17 20 gnd NMOS_VTL L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06 $X=6325 $Y=600 $D=1
M13 21 R gnd gnd NMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06 $X=6785 $Y=600 $D=1
M14 17 16 21 gnd NMOS_VTL L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06 $X=7165 $Y=600 $D=1
M15 Q 17 gnd gnd NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07 $X=7970 $Y=355 $D=1
M16 vdd CLK 10 8 PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06 $X=635 $Y=2370 $D=0
M17 11 D vdd 8 PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06 $X=1165 $Y=2370 $D=0
M18 13 9 11 8 PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14 PD=1.09e-06 PS=1.28e-06 $X=1545 $Y=2370 $D=0
M19 12 10 13 8 PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14 PD=1.38e-06 PS=1.09e-06 $X=2235 $Y=2370 $D=0
M20 vdd 10 9 8 PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06 $X=2235 $Y=3585 $D=0
M21 vdd R 12 8 PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06 $X=2715 $Y=2370 $D=0
M22 12 14 vdd 8 PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13 PD=1.21e-06 PS=2.33e-06 $X=3275 $Y=2370 $D=0
M23 14 S vdd 8 PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06 $X=4315 $Y=2625 $D=0
M24 16 10 14 8 PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13 PD=7.8e-07 PS=3.12e-06 $X=5065 $Y=2625 $D=0
M25 vdd 13 14 8 PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06 PS=3.12e-06 $X=5065 $Y=3495 $D=0
M26 15 9 16 8 PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14 PD=3.3e-06 PS=7.8e-07 $X=5445 $Y=2625 $D=0
M27 15 17 vdd 8 PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06 PS=1.28e-06 $X=5445 $Y=3495 $D=0
M28 vdd S 15 8 PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06 $X=6305 $Y=2625 $D=0
M29 17 R vdd 8 PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06 $X=6785 $Y=2625 $D=0
M30 vdd 16 17 8 PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06 PS=1.28e-06 $X=7165 $Y=2625 $D=0
M31 Q 17 vdd 8 PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06 $X=7675 $Y=2625 $D=0
.ENDS
***************************************
.SUBCKT fullsystem
** N=49 EP=0 IP=309 FDC=322
M0 45 12 32 32 NMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.21e-06 $X=60560 $Y=55455 $D=1
M1 20 13 45 32 NMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=7e-14 PD=1.28e-06 PS=1.28e-06 $X=60940 $Y=55455 $D=1
M2 46 14 20 32 NMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=7e-14 PD=1.28e-06 PS=1.28e-06 $X=61320 $Y=55455 $D=1
M3 32 21 46 32 NMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06 $X=61700 $Y=55455 $D=1
M4 47 28 31 32 NMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.21e-06 $X=62655 $Y=55495 $D=1
M5 32 16 47 32 NMOS_VTL L=5e-08 W=5e-07 AD=1.175e-13 AS=7e-14 PD=1.47e-06 PS=1.28e-06 $X=63035 $Y=55495 $D=1
M6 32 21 33 32 NMOS_VTL L=5e-08 W=5e-07 AD=1.225e-13 AS=5.25e-14 PD=1.515e-06 PS=1.21e-06 $X=63385 $Y=65660 $D=1
M7 17 31 32 32 NMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.175e-13 PD=1.21e-06 PS=1.47e-06 $X=63605 $Y=55495 $D=1
M8 48 21 32 32 NMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.225e-13 PD=1.28e-06 PS=1.515e-06 $X=63975 $Y=65635 $D=1
M9 16 19 48 32 NMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=7e-14 PD=1.28e-06 PS=1.28e-06 $X=64355 $Y=65635 $D=1
M10 49 36 16 32 NMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=7e-14 PD=1.28e-06 PS=1.28e-06 $X=64735 $Y=65635 $D=1
M11 32 33 49 32 NMOS_VTL L=5e-08 W=5e-07 AD=2.025e-13 AS=7e-14 PD=1.81e-06 PS=1.28e-06 $X=65115 $Y=65635 $D=1
M12 34 19 32 32 NMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=2.625e-14 PD=7.8e-07 PS=7.1e-07 $X=65120 $Y=46075 $D=1
M13 32 20 34 32 NMOS_VTL L=5e-08 W=2.5e-07 AD=7.875e-14 AS=3.5e-14 PD=1.49e-06 PS=7.8e-07 $X=65500 $Y=46075 $D=1
M14 36 19 32 32 NMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=2.025e-13 PD=1.21e-06 PS=1.81e-06 $X=66025 $Y=65635 $D=1
M15 37 34 32 32 NMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=7.875e-14 PD=1.21e-06 PS=1.49e-06 $X=66090 $Y=45575 $D=1
M16 38 21 32 32 NMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=2.625e-14 PD=7.8e-07 PS=7.1e-07 $X=67400 $Y=65335 $D=1
M17 32 16 38 32 NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=3.5e-14 PD=7.1e-07 PS=7.8e-07 $X=67780 $Y=65335 $D=1
M18 20 12 30 22 PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13 AS=1.05e-13 PD=2.28e-06 PS=2.21e-06 $X=60560 $Y=57345 $D=0
M19 30 13 20 22 PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13 AS=1.4e-13 PD=2.28e-06 PS=2.28e-06 $X=60940 $Y=57345 $D=0
M20 22 14 30 22 PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13 AS=1.4e-13 PD=2.28e-06 PS=2.28e-06 $X=61320 $Y=57345 $D=0
M21 30 21 22 22 PMOS_VTL L=5e-08 W=1e-06 AD=1.05e-13 AS=1.4e-13 PD=2.21e-06 PS=2.28e-06 $X=61700 $Y=57345 $D=0
M22 31 28 22 22 PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.21e-06 $X=62655 $Y=57680 $D=0
M23 22 16 31 22 PMOS_VTL L=5e-08 W=5e-07 AD=1.575e-13 AS=7e-14 PD=2.49e-06 PS=1.28e-06 $X=63035 $Y=57680 $D=0
M24 22 21 33 22 PMOS_VTL L=5e-08 W=1e-06 AD=3.05e-13 AS=1.05e-13 PD=2.61e-06 PS=2.21e-06 $X=63385 $Y=67565 $D=0
M25 17 31 22 22 PMOS_VTL L=5e-08 W=1e-06 AD=1.05e-13 AS=1.575e-13 PD=2.21e-06 PS=2.49e-06 $X=63625 $Y=57680 $D=0
M26 41 21 22 22 PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13 AS=3.05e-13 PD=2.28e-06 PS=2.61e-06 $X=64095 $Y=67565 $D=0
M27 16 36 41 22 PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13 AS=1.4e-13 PD=2.28e-06 PS=2.28e-06 $X=64475 $Y=67565 $D=0
M28 42 19 16 22 PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13 AS=1.4e-13 PD=2.28e-06 PS=2.28e-06 $X=64855 $Y=67565 $D=0
M29 43 19 34 22 PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13 AS=1.05e-13 PD=2.28e-06 PS=2.21e-06 $X=65120 $Y=47800 $D=0
M30 22 33 42 22 PMOS_VTL L=5e-08 W=1e-06 AD=3.45e-13 AS=1.4e-13 PD=2.69e-06 PS=2.28e-06 $X=65235 $Y=67565 $D=0
M31 22 20 43 22 PMOS_VTL L=5e-08 W=1e-06 AD=2.45e-13 AS=1.4e-13 PD=2.49e-06 PS=2.28e-06 $X=65500 $Y=47800 $D=0
M32 36 19 22 22 PMOS_VTL L=5e-08 W=1e-06 AD=1.05e-13 AS=3.45e-13 PD=2.21e-06 PS=2.69e-06 $X=66025 $Y=67565 $D=0
M33 37 34 22 22 PMOS_VTL L=5e-08 W=1e-06 AD=1.05e-13 AS=2.45e-13 PD=2.21e-06 PS=2.49e-06 $X=66090 $Y=47800 $D=0
M34 44 21 22 22 PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13 AS=1.05e-13 PD=2.28e-06 PS=2.21e-06 $X=67400 $Y=66325 $D=0
M35 38 16 44 22 PMOS_VTL L=5e-08 W=1e-06 AD=1.05e-13 AS=1.4e-13 PD=2.21e-06 PS=2.28e-06 $X=67780 $Y=66325 $D=0
X188 23 32 22 2 INVX1 $T=42560 64980 0 0 $X=42360 $Y=64780
X189 7 32 22 24 INVX1 $T=45600 55100 1 0 $X=45400 $Y=49960
X190 25 32 22 3 INVX1 $T=48640 64980 0 0 $X=48440 $Y=64780
X191 6 32 22 25 INVX1 $T=50160 64980 0 0 $X=49960 $Y=64780
X192 9 32 22 26 INVX1 $T=51680 45220 1 0 $X=51480 $Y=40080
X193 28 32 22 14 INVX1 $T=60800 55100 1 0 $X=60600 $Y=49960
X194 32 22 15 23 ICV_4 $T=40280 64980 0 0 $X=40080 $Y=64780
X195 32 22 24 5 ICV_4 $T=43320 55100 1 0 $X=43120 $Y=49960
X196 32 22 26 8 ICV_4 $T=49400 45220 1 0 $X=49200 $Y=40080
X197 32 22 27 10 ICV_4 $T=53960 45220 0 0 $X=53760 $Y=45020
X198 32 22 21 13 ICV_4 $T=56240 55100 0 0 $X=56040 $Y=54900
X199 32 22 18 27 ICV_4 $T=57760 45220 1 0 $X=57560 $Y=40080
X200 32 22 39 29 ICV_4 $T=57760 64980 0 0 $X=57560 $Y=64780
X201 32 22 40 35 ICV_4 $T=64600 55100 0 0 $X=64400 $Y=54900
X202 32 22 37 11 ICV_4 $T=66880 45220 0 0 $X=66680 $Y=45020
X203 1 2 22 29 22 32 6 22 DFFSR $T=42560 64980 1 0 $X=42360 $Y=59840
X204 1 3 22 29 22 32 7 22 DFFSR $T=43320 55100 0 0 $X=43120 $Y=54900
X205 4 5 22 35 22 32 9 22 DFFSR $T=44080 45220 0 0 $X=43880 $Y=45020
X206 4 8 22 35 22 32 28 22 DFFSR $T=50920 55100 1 0 $X=50720 $Y=49960
X207 1 10 22 29 22 32 15 22 DFFSR $T=53960 64980 1 0 $X=53760 $Y=59840
X208 4 11 22 35 22 32 18 22 DFFSR $T=56240 45220 0 0 $X=56040 $Y=45020
X209 4 11 22 35 22 32 21 22 DFFSR $T=62320 55100 1 0 $X=62120 $Y=49960
X210 4 17 22 35 22 32 19 22 DFFSR $T=62320 64980 1 0 $X=62120 $Y=59840
.ENDS
***************************************
