* File: /media/ntfsdrive1/workspace/ProjectDIC2/runsets/pex/extracted.sp
* Created: Mon Dec  7 09:37:15 2015
* Program "Calibre xRC"
* Version "v2013.3_28.19"
* 
.include "/media/ntfsdrive1/workspace/ProjectDIC2/runsets/pex/extracted.sp.pex"
.subckt FULLSYSTEM 
* 
M0 N_17_M0_d N_4_M0_g N_1_M0_s N_1_X153/M0_b NMOS_VTL L=5e-08 W=2.5e-07
+ AD=3.5e-14 AS=2.625e-14 PD=7.8e-07 PS=7.1e-07
M1 N_1_M1_d N_7_M1_g N_17_M0_d N_1_X153/M0_b NMOS_VTL L=5e-08 W=2.5e-07
+ AD=2.625e-14 AS=3.5e-14 PD=7.1e-07 PS=7.8e-07
M2 N_1_M2_s N_21_M2_g N_1_M2_s N_1_X153/M0_b NMOS_VTL L=5e-08 W=5e-07
+ AD=1.225e-13 AS=5.25e-14 PD=1.515e-06 PS=1.21e-06
M3 46 N_20_M3_g N_7_M3_s N_1_X156/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=7e-14
+ AS=5.25e-14 PD=1.28e-06 PS=1.21e-06
M4 N_1_M4_s N_18_M4_g N_1_M4_s N_1_X154/M0_b NMOS_VTL L=5e-08 W=2.5e-07
+ AD=3.5e-14 AS=2.625e-14 PD=7.8e-07 PS=7.1e-07
M5 47 N_19_M5_g N_1_M5_s N_1_X156/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=7e-14
+ AS=5.25e-14 PD=1.28e-06 PS=1.21e-06
M6 N_1_M6_d N_22_M6_g 46 N_1_X156/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=1.175e-13
+ AS=7e-14 PD=1.47e-06 PS=1.28e-06
M7 48 N_21_M7_g N_1_M2_s N_1_X153/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=7e-14
+ AS=1.225e-13 PD=1.28e-06 PS=1.515e-06
M8 N_1_M4_s N_1_M8_g N_1_M4_s N_1_X154/M0_b NMOS_VTL L=5e-08 W=2.5e-07
+ AD=7.875e-14 AS=3.5e-14 PD=1.49e-06 PS=7.8e-07
M9 N_23_M9_d N_8_M9_g 47 N_1_X156/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=7e-14
+ AS=7e-14 PD=1.28e-06 PS=1.28e-06
M10 N_24_M10_d N_7_M10_g 48 N_1_X153/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=7e-14
+ AS=7e-14 PD=1.28e-06 PS=1.28e-06
M11 49 N_9_M11_g N_23_M9_d N_1_X156/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=7e-14
+ AS=7e-14 PD=1.28e-06 PS=1.28e-06
M12 N_25_M12_d N_7_M12_g N_1_M6_d N_1_X156/M0_b NMOS_VTL L=5e-08 W=5e-07
+ AD=5.25e-14 AS=1.175e-13 PD=1.21e-06 PS=1.47e-06
M13 N_1_M4_s N_1_M13_g N_1_M4_s N_1_X154/M0_b NMOS_VTL L=5e-08 W=5e-07
+ AD=5.25e-14 AS=7.875e-14 PD=1.21e-06 PS=1.49e-06
M14 50 N_27_M14_g N_24_M10_d N_1_X153/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=7e-14
+ AS=7e-14 PD=1.28e-06 PS=1.28e-06
M15 N_1_M15_d N_4_M15_g 49 N_1_X156/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14
+ AS=7e-14 PD=1.21e-06 PS=1.28e-06
M16 N_1_M16_d N_1_M16_g 50 N_1_X153/M0_b NMOS_VTL L=5e-08 W=5e-07 AD=2.025e-13
+ AS=7e-14 PD=1.81e-06 PS=1.28e-06
M17 N_27_M17_d N_7_M17_g N_1_M16_d N_1_X153/M0_b NMOS_VTL L=5e-08 W=5e-07
+ AD=5.25e-14 AS=2.025e-13 PD=1.21e-06 PS=1.81e-06
M18 N_1_M18_s N_1_M18_g N_1_M18_s N_1_X153/M0_b NMOS_VTL L=5e-08 W=5e-07
+ AD=8.75e-14 AS=5.25e-14 PD=1.49e-06 PS=1.21e-06
M19 N_1_M18_s N_1_M19_g N_1_M18_s N_1_X153/M0_b NMOS_VTL L=5e-08 W=2.5e-07
+ AD=2.625e-14 AS=8.75e-14 PD=7.1e-07 PS=1.49e-06
M20 N_6_M20_d N_28_M20_g N_1_M20_s N_1_X153/M0_b NMOS_VTL L=5e-08 W=5e-07
+ AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
M21 42 N_4_M21_g N_5_M21_s N_5_X156/M16_b PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13
+ AS=1.05e-13 PD=2.28e-06 PS=2.21e-06
M22 N_17_M22_d N_7_M22_g 42 N_5_X156/M16_b PMOS_VTL L=5e-08 W=1e-06 AD=1.05e-13
+ AS=1.4e-13 PD=2.21e-06 PS=2.28e-06
M23 N_5_M23_d N_21_M23_g N_1_M23_s N_5_X153/M16_b PMOS_VTL L=5e-08 W=1e-06
+ AD=3.05e-13 AS=1.05e-13 PD=2.61e-06 PS=2.21e-06
M24 N_7_M24_d N_20_M24_g N_5_M24_s N_5_X156/M16_b PMOS_VTL L=5e-08 W=5e-07
+ AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.21e-06
M25 43 N_18_M25_g N_1_M25_s N_5_X158/M16_b PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13
+ AS=1.05e-13 PD=2.28e-06 PS=2.21e-06
M26 N_23_M26_d N_19_M26_g N_26_M26_s N_5_X162/M3_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.4e-13 AS=1.05e-13 PD=2.28e-06 PS=2.21e-06
M27 N_5_M27_d N_22_M27_g N_7_M24_d N_5_X156/M16_b PMOS_VTL L=5e-08 W=5e-07
+ AD=1.575e-13 AS=7e-14 PD=2.49e-06 PS=1.28e-06
M28 N_5_M28_d N_1_M28_g 43 N_5_X158/M16_b PMOS_VTL L=5e-08 W=1e-06 AD=2.45e-13
+ AS=1.4e-13 PD=2.49e-06 PS=2.28e-06
M29 N_26_M29_d N_8_M29_g N_23_M26_d N_5_X162/M3_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.4e-13 AS=1.4e-13 PD=2.28e-06 PS=2.28e-06
M30 44 N_21_M30_g N_5_M23_d N_5_X153/M16_b PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13
+ AS=3.05e-13 PD=2.28e-06 PS=2.61e-06
M31 N_5_M31_d N_9_M31_g N_26_M29_d N_5_X162/M3_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.4e-13 AS=1.4e-13 PD=2.28e-06 PS=2.28e-06
M32 N_25_M32_d N_7_M32_g N_5_M27_d N_5_X156/M16_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.05e-13 AS=1.575e-13 PD=2.21e-06 PS=2.49e-06
M33 N_24_M33_d N_27_M33_g 44 N_5_X153/M16_b PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13
+ AS=1.4e-13 PD=2.28e-06 PS=2.28e-06
M34 N_1_M34_d N_1_M34_g N_5_M28_d N_5_X158/M16_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.05e-13 AS=2.45e-13 PD=2.21e-06 PS=2.49e-06
M35 N_26_M35_d N_4_M35_g N_5_M31_d N_5_X162/M3_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.05e-13 AS=1.4e-13 PD=2.21e-06 PS=2.28e-06
M36 45 N_7_M36_g N_24_M33_d N_5_X153/M16_b PMOS_VTL L=5e-08 W=1e-06 AD=1.4e-13
+ AS=1.4e-13 PD=2.28e-06 PS=2.28e-06
M37 N_5_M37_d N_1_M37_g 45 N_5_X153/M16_b PMOS_VTL L=5e-08 W=1e-06 AD=3.45e-13
+ AS=1.4e-13 PD=2.69e-06 PS=2.28e-06
M38 N_27_M38_d N_7_M38_g N_5_M37_d N_5_X153/M16_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.05e-13 AS=3.45e-13 PD=2.21e-06 PS=2.69e-06
M39 N_5_M39_d N_1_M39_g N_1_M39_s N_5_X153/M16_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.75e-13 AS=1.05e-13 PD=2.49e-06 PS=2.21e-06
M40 N_1_M40_d N_1_M40_g N_5_M39_d N_5_X153/M16_b PMOS_VTL L=5e-08 W=5e-07
+ AD=5.25e-14 AS=1.75e-13 PD=1.21e-06 PS=2.49e-06
M41 N_6_M41_d N_28_M41_g N_5_M41_s N_5_X156/M16_b PMOS_VTL L=5e-08 W=1e-06
+ AD=1.05e-13 AS=1.05e-13 PD=2.21e-06 PS=2.21e-06
mX153/M0 N_1_X153/M0_s N_X153/CLK_X153/M0_g N_1_X153/M0_s N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX153/M1 N_X153/11_X153/M1_d N_X153/D_X153/M1_g N_1_X153/M0_s N_1_X153/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX153/M2 N_29_X153/M2_d N_1_X153/M2_g N_1_X153/M2_s N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX153/M3 N_X153/13_X153/M3_d N_1_X153/M3_g N_X153/11_X153/M1_d N_1_X153/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06 PS=9.2e-07
mX153/M4 N_X153/12_X153/M4_d N_29_X153/M4_g N_X153/13_X153/M3_d N_1_X153/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06 PS=1.2e-06
mX153/M5 X153/17 N_6_X153/M5_g N_X153/12_X153/M4_d N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX153/M6 N_1_X153/M6_d N_X153/14_X153/M6_g X153/17 N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX153/M7 X153/18 N_X153/13_X153/M7_g N_1_X153/M6_d N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX153/M8 N_X153/14_X153/M8_d N_5_X153/M8_g X153/18 N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX153/M9 N_1_X153/M9_d N_29_X153/M9_g N_X153/14_X153/M8_d N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06 PS=1.38e-06
mX153/M10 N_X153/15_X153/M10_d N_1_X153/M10_g N_1_X153/M9_d N_1_X153/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06 PS=1.04e-06
mX153/M11 X153/19 N_5_X153/M11_g N_X153/15_X153/M10_d N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX153/M12 N_1_X153/M12_d N_X153/16_X153/M12_g X153/19 N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX153/M13 X153/20 N_6_X153/M13_g N_1_X153/M12_d N_1_X153/M0_b NMOS_VTL L=5e-08
+ W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX153/M14 N_X153/16_X153/M14_d N_1_X153/M14_g X153/20 N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX153/M15 N_4_X153/M15_d N_X153/16_X153/M15_g N_1_X153/M15_s N_1_X153/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX153/M16 N_5_X153/M16_d N_X153/CLK_X153/M16_g N_1_X153/M16_s N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX153/M17 N_X153/11_X153/M17_d N_X153/D_X153/M17_g N_5_X153/M16_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX153/M18 N_X153/13_X153/M18_d N_29_X153/M18_g N_X153/11_X153/M17_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14 PD=1.09e-06
+ PS=1.28e-06
mX153/M19 N_X153/12_X153/M19_d N_1_X153/M19_g N_X153/13_X153/M18_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14 PD=1.38e-06
+ PS=1.09e-06
mX153/M20 N_5_X153/M20_d N_1_X153/M20_g N_29_X153/M20_s N_5_X153/M16_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX153/M21 N_5_X153/M21_d N_6_X153/M21_g N_X153/12_X153/M19_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX153/M22 N_X153/12_X153/M22_d N_X153/14_X153/M22_g N_5_X153/M21_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13 PD=1.21e-06
+ PS=2.33e-06
mX153/M23 N_X153/14_X153/M23_d N_5_X153/M23_g N_5_X153/M23_s N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX153/M24 N_1_X153/M24_d N_1_X153/M24_g N_X153/14_X153/M23_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13 PD=7.8e-07 PS=3.12e-06
mX153/M25 N_5_X153/M25_d N_X153/13_X153/M25_g N_X153/14_X153/M23_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX153/M26 N_X153/15_X153/M26_d N_29_X153/M26_g N_1_X153/M24_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14 PD=3.3e-06 PS=7.8e-07
mX153/M27 N_X153/15_X153/M26_d N_X153/16_X153/M27_g N_5_X153/M25_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX153/M28 N_5_X153/M28_d N_5_X153/M28_g N_X153/15_X153/M26_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX153/M29 N_X153/16_X153/M29_d N_6_X153/M29_g N_5_X153/M28_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX153/M30 N_5_X153/M30_d N_1_X153/M30_g N_X153/16_X153/M29_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06 PS=1.28e-06
mX153/M31 N_4_X153/M31_d N_X153/16_X153/M31_g N_5_X153/M30_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
mX154/M0 N_1_X154/M0_s N_X154/CLK_X154/M0_g N_1_X154/M0_s N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX154/M1 N_X154/11_X154/M1_d N_X154/D_X154/M1_g N_1_X154/M0_s N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX154/M2 N_5_X154/M2_d N_1_X154/M2_g N_1_X154/M2_s N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX154/M3 N_X154/13_X154/M3_d N_1_X154/M3_g N_X154/11_X154/M1_d N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06 PS=9.2e-07
mX154/M4 N_X154/12_X154/M4_d N_5_X154/M4_g N_X154/13_X154/M3_d N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06 PS=1.2e-06
mX154/M5 X154/17 N_6_X154/M5_g N_X154/12_X154/M4_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX154/M6 N_1_X154/M6_d N_X154/14_X154/M6_g X154/17 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX154/M7 X154/18 N_X154/13_X154/M7_g N_1_X154/M6_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX154/M8 N_X154/14_X154/M8_d N_5_X154/M8_g X154/18 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX154/M9 N_30_X154/M9_d N_5_X154/M9_g N_X154/14_X154/M8_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06 PS=1.38e-06
mX154/M10 N_X154/15_X154/M10_d N_1_X154/M10_g N_30_X154/M9_d N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06 PS=1.04e-06
mX154/M11 X154/19 N_5_X154/M11_g N_X154/15_X154/M10_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX154/M12 N_1_X154/M12_d N_X154/16_X154/M12_g X154/19 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX154/M13 X154/20 N_6_X154/M13_g N_1_X154/M12_d N_1_X154/M0_b NMOS_VTL L=5e-08
+ W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX154/M14 N_X154/16_X154/M14_d N_30_X154/M14_g X154/20 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX154/M15 N_11_X154/M15_d N_X154/16_X154/M15_g N_1_X154/M15_s N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX154/M16 N_5_X154/M16_d N_X154/CLK_X154/M16_g N_1_X154/M16_s N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX154/M17 N_X154/11_X154/M17_d N_X154/D_X154/M17_g N_5_X154/M16_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX154/M18 N_X154/13_X154/M18_d N_5_X154/M18_g N_X154/11_X154/M17_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14 PD=1.09e-06
+ PS=1.28e-06
mX154/M19 N_X154/12_X154/M19_d N_1_X154/M19_g N_X154/13_X154/M18_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14 PD=1.38e-06
+ PS=1.09e-06
mX154/M20 N_5_X154/M20_d N_1_X154/M20_g N_5_X154/M20_s N_5_X153/M16_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX154/M21 N_5_X154/M21_d N_6_X154/M21_g N_X154/12_X154/M19_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX154/M22 N_X154/12_X154/M22_d N_X154/14_X154/M22_g N_5_X154/M21_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13 PD=1.21e-06
+ PS=2.33e-06
mX154/M23 N_X154/14_X154/M23_d N_5_X154/M23_g N_5_X154/M23_s N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX154/M24 N_30_X154/M24_d N_1_X154/M24_g N_X154/14_X154/M23_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13 PD=7.8e-07 PS=3.12e-06
mX154/M25 N_5_X154/M25_d N_X154/13_X154/M25_g N_X154/14_X154/M23_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX154/M26 N_X154/15_X154/M26_d N_5_X154/M26_g N_30_X154/M24_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14 PD=3.3e-06 PS=7.8e-07
mX154/M27 N_X154/15_X154/M26_d N_X154/16_X154/M27_g N_5_X154/M25_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX154/M28 N_5_X154/M28_d N_5_X154/M28_g N_X154/15_X154/M26_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX154/M29 N_X154/16_X154/M29_d N_6_X154/M29_g N_5_X154/M28_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX154/M30 N_5_X154/M30_d N_30_X154/M30_g N_X154/16_X154/M29_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06 PS=1.28e-06
mX154/M31 N_11_X154/M31_d N_X154/16_X154/M31_g N_5_X154/M30_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
mX155/M0 N_1_X155/M0_s N_X155/CLK_X155/M0_g N_1_X155/M0_s N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX155/M1 N_X155/11_X155/M1_d N_X155/D_X155/M1_g N_1_X155/M0_s N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX155/M2 N_5_X155/M2_d N_1_X155/M2_g N_1_X155/M2_s N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX155/M3 N_X155/13_X155/M3_d N_1_X155/M3_g N_X155/11_X155/M1_d N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06 PS=9.2e-07
mX155/M4 N_X155/12_X155/M4_d N_5_X155/M4_g N_X155/13_X155/M3_d N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06 PS=1.2e-06
mX155/M5 X155/17 N_6_X155/M5_g N_X155/12_X155/M4_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX155/M6 N_1_X155/M6_d N_X155/14_X155/M6_g X155/17 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX155/M7 X155/18 N_X155/13_X155/M7_g N_1_X155/M6_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX155/M8 N_X155/14_X155/M8_d N_5_X155/M8_g X155/18 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX155/M9 N_31_X155/M9_d N_5_X155/M9_g N_X155/14_X155/M8_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06 PS=1.38e-06
mX155/M10 N_X155/15_X155/M10_d N_1_X155/M10_g N_31_X155/M9_d N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06 PS=1.04e-06
mX155/M11 X155/19 N_5_X155/M11_g N_X155/15_X155/M10_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX155/M12 N_1_X155/M12_d N_X155/16_X155/M12_g X155/19 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX155/M13 X155/20 N_6_X155/M13_g N_1_X155/M12_d N_1_X154/M0_b NMOS_VTL L=5e-08
+ W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX155/M14 N_X155/16_X155/M14_d N_31_X155/M14_g X155/20 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX155/M15 N_7_X155/M15_d N_X155/16_X155/M15_g N_1_X155/M15_s N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX155/M16 N_5_X155/M16_d N_X155/CLK_X155/M16_g N_1_X155/M16_s N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX155/M17 N_X155/11_X155/M17_d N_X155/D_X155/M17_g N_5_X155/M16_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX155/M18 N_X155/13_X155/M18_d N_5_X155/M18_g N_X155/11_X155/M17_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14 PD=1.09e-06
+ PS=1.28e-06
mX155/M19 N_X155/12_X155/M19_d N_1_X155/M19_g N_X155/13_X155/M18_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14 PD=1.38e-06
+ PS=1.09e-06
mX155/M20 N_5_X155/M20_d N_1_X155/M20_g N_5_X155/M20_s N_5_X153/M16_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX155/M21 N_5_X155/M21_d N_6_X155/M21_g N_X155/12_X155/M19_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX155/M22 N_X155/12_X155/M22_d N_X155/14_X155/M22_g N_5_X155/M21_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13 PD=1.21e-06
+ PS=2.33e-06
mX155/M23 N_X155/14_X155/M23_d N_5_X155/M23_g N_5_X155/M23_s N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX155/M24 N_31_X155/M24_d N_1_X155/M24_g N_X155/14_X155/M23_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13 PD=7.8e-07 PS=3.12e-06
mX155/M25 N_5_X155/M25_d N_X155/13_X155/M25_g N_X155/14_X155/M23_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX155/M26 N_X155/15_X155/M26_d N_5_X155/M26_g N_31_X155/M24_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14 PD=3.3e-06 PS=7.8e-07
mX155/M27 N_X155/15_X155/M26_d N_X155/16_X155/M27_g N_5_X155/M25_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX155/M28 N_5_X155/M28_d N_5_X155/M28_g N_X155/15_X155/M26_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX155/M29 N_X155/16_X155/M29_d N_6_X155/M29_g N_5_X155/M28_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX155/M30 N_5_X155/M30_d N_31_X155/M30_g N_X155/16_X155/M29_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06 PS=1.28e-06
mX155/M31 N_7_X155/M31_d N_X155/16_X155/M31_g N_5_X155/M30_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
mX156/M0 N_1_X156/M0_s N_X156/CLK_X156/M0_g N_1_X156/M0_s N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX156/M1 N_X156/11_X156/M1_d N_X156/D_X156/M1_g N_1_X156/M0_s N_1_X156/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX156/M2 N_32_X156/M2_d N_1_X156/M2_g N_1_X156/M2_s N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX156/M3 N_X156/13_X156/M3_d N_1_X156/M3_g N_X156/11_X156/M1_d N_1_X156/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06 PS=9.2e-07
mX156/M4 N_X156/12_X156/M4_d N_32_X156/M4_g N_X156/13_X156/M3_d N_1_X156/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06 PS=1.2e-06
mX156/M5 X156/17 N_14_X156/M5_g N_X156/12_X156/M4_d N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX156/M6 N_1_X156/M6_d N_X156/14_X156/M6_g X156/17 N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX156/M7 X156/18 N_X156/13_X156/M7_g N_1_X156/M6_d N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX156/M8 N_X156/14_X156/M8_d N_5_X156/M8_g X156/18 N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX156/M9 N_1_X156/M9_d N_32_X156/M9_g N_X156/14_X156/M8_d N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06 PS=1.38e-06
mX156/M10 N_X156/15_X156/M10_d N_1_X156/M10_g N_1_X156/M9_d N_1_X156/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06 PS=1.04e-06
mX156/M11 X156/19 N_5_X156/M11_g N_X156/15_X156/M10_d N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX156/M12 N_1_X156/M12_d N_X156/16_X156/M12_g X156/19 N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX156/M13 X156/20 N_14_X156/M13_g N_1_X156/M12_d N_1_X156/M0_b NMOS_VTL L=5e-08
+ W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX156/M14 N_X156/16_X156/M14_d N_1_X156/M14_g X156/20 N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX156/M15 N_1_X156/M15_d N_X156/16_X156/M15_g N_1_X156/M15_s N_1_X156/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX156/M16 N_5_X156/M16_d N_X156/CLK_X156/M16_g N_1_X156/M16_s N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX156/M17 N_X156/11_X156/M17_d N_X156/D_X156/M17_g N_5_X156/M16_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX156/M18 N_X156/13_X156/M18_d N_32_X156/M18_g N_X156/11_X156/M17_d
+ N_5_X156/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14 PD=1.09e-06
+ PS=1.28e-06
mX156/M19 N_X156/12_X156/M19_d N_1_X156/M19_g N_X156/13_X156/M18_d
+ N_5_X156/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14 PD=1.38e-06
+ PS=1.09e-06
mX156/M20 N_5_X156/M20_d N_1_X156/M20_g N_32_X156/M20_s N_5_X156/M16_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX156/M21 N_5_X156/M21_d N_14_X156/M21_g N_X156/12_X156/M19_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX156/M22 N_X156/12_X156/M22_d N_X156/14_X156/M22_g N_5_X156/M21_d
+ N_5_X156/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13 PD=1.21e-06
+ PS=2.33e-06
mX156/M23 N_X156/14_X156/M23_d N_5_X156/M23_g N_5_X156/M23_s N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX156/M24 N_1_X156/M24_d N_1_X156/M24_g N_X156/14_X156/M23_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13 PD=7.8e-07 PS=3.12e-06
mX156/M25 N_5_X156/M25_d N_X156/13_X156/M25_g N_X156/14_X156/M23_d
+ N_5_X156/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX156/M26 N_X156/15_X156/M26_d N_32_X156/M26_g N_1_X156/M24_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14 PD=3.3e-06 PS=7.8e-07
mX156/M27 N_X156/15_X156/M26_d N_X156/16_X156/M27_g N_5_X156/M25_d
+ N_5_X156/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX156/M28 N_5_X156/M28_d N_5_X156/M28_g N_X156/15_X156/M26_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX156/M29 N_X156/16_X156/M29_d N_14_X156/M29_g N_5_X156/M28_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX156/M30 N_5_X156/M30_d N_1_X156/M30_g N_X156/16_X156/M29_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06 PS=1.28e-06
mX156/M31 N_1_X156/M31_d N_X156/16_X156/M31_g N_5_X156/M30_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
mX157/M0 N_1_X157/M0_s N_X157/CLK_X157/M0_g N_1_X157/M0_s N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX157/M1 N_X157/11_X157/M1_d N_X157/D_X157/M1_g N_1_X157/M0_s N_1_X153/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX157/M2 N_5_X157/M2_d N_1_X157/M2_g N_1_X157/M2_s N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX157/M3 N_X157/13_X157/M3_d N_1_X157/M3_g N_X157/11_X157/M1_d N_1_X153/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06 PS=9.2e-07
mX157/M4 N_X157/12_X157/M4_d N_5_X157/M4_g N_X157/13_X157/M3_d N_1_X153/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06 PS=1.2e-06
mX157/M5 X157/17 N_14_X157/M5_g N_X157/12_X157/M4_d N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX157/M6 N_1_X157/M6_d N_X157/14_X157/M6_g X157/17 N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX157/M7 X157/18 N_X157/13_X157/M7_g N_1_X157/M6_d N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX157/M8 N_X157/14_X157/M8_d N_5_X157/M8_g X157/18 N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX157/M9 N_33_X157/M9_d N_5_X157/M9_g N_X157/14_X157/M8_d N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06 PS=1.38e-06
mX157/M10 N_X157/15_X157/M10_d N_1_X157/M10_g N_33_X157/M9_d N_1_X153/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06 PS=1.04e-06
mX157/M11 X157/19 N_5_X157/M11_g N_X157/15_X157/M10_d N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX157/M12 N_1_X157/M12_d N_X157/16_X157/M12_g X157/19 N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX157/M13 X157/20 N_14_X157/M13_g N_1_X157/M12_d N_1_X153/M0_b NMOS_VTL L=5e-08
+ W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX157/M14 N_X157/16_X157/M14_d N_33_X157/M14_g X157/20 N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX157/M15 N_34_X157/M15_d N_X157/16_X157/M15_g N_1_X157/M15_s N_1_X153/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX157/M16 N_5_X157/M16_d N_X157/CLK_X157/M16_g N_1_X157/M16_s N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX157/M17 N_X157/11_X157/M17_d N_X157/D_X157/M17_g N_5_X157/M16_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX157/M18 N_X157/13_X157/M18_d N_5_X157/M18_g N_X157/11_X157/M17_d
+ N_5_X156/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14 PD=1.09e-06
+ PS=1.28e-06
mX157/M19 N_X157/12_X157/M19_d N_1_X157/M19_g N_X157/13_X157/M18_d
+ N_5_X156/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14 PD=1.38e-06
+ PS=1.09e-06
mX157/M20 N_5_X157/M20_d N_1_X157/M20_g N_5_X157/M20_s N_5_X156/M16_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX157/M21 N_5_X157/M21_d N_14_X157/M21_g N_X157/12_X157/M19_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX157/M22 N_X157/12_X157/M22_d N_X157/14_X157/M22_g N_5_X157/M21_d
+ N_5_X156/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13 PD=1.21e-06
+ PS=2.33e-06
mX157/M23 N_X157/14_X157/M23_d N_5_X157/M23_g N_5_X157/M23_s N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX157/M24 N_33_X157/M24_d N_1_X157/M24_g N_X157/14_X157/M23_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13 PD=7.8e-07 PS=3.12e-06
mX157/M25 N_5_X157/M25_d N_X157/13_X157/M25_g N_X157/14_X157/M23_d
+ N_5_X156/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX157/M26 N_X157/15_X157/M26_d N_5_X157/M26_g N_33_X157/M24_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14 PD=3.3e-06 PS=7.8e-07
mX157/M27 N_X157/15_X157/M26_d N_X157/16_X157/M27_g N_5_X157/M25_d
+ N_5_X156/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX157/M28 N_5_X157/M28_d N_5_X157/M28_g N_X157/15_X157/M26_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX157/M29 N_X157/16_X157/M29_d N_14_X157/M29_g N_5_X157/M28_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX157/M30 N_5_X157/M30_d N_33_X157/M30_g N_X157/16_X157/M29_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06 PS=1.28e-06
mX157/M31 N_34_X157/M31_d N_X157/16_X157/M31_g N_5_X157/M30_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
mX158/M0 N_1_X158/M0_s N_X158/CLK_X158/M0_g N_1_X158/M0_s N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX158/M1 N_X158/11_X158/M1_d N_X158/D_X158/M1_g N_1_X158/M0_s N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX158/M2 N_35_X158/M2_d N_1_X158/M2_g N_1_X158/M2_s N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX158/M3 N_X158/13_X158/M3_d N_1_X158/M3_g N_X158/11_X158/M1_d N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06 PS=9.2e-07
mX158/M4 N_X158/12_X158/M4_d N_35_X158/M4_g N_X158/13_X158/M3_d N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06 PS=1.2e-06
mX158/M5 X158/17 N_6_X158/M5_g N_X158/12_X158/M4_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX158/M6 N_1_X158/M6_d N_X158/14_X158/M6_g X158/17 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX158/M7 X158/18 N_X158/13_X158/M7_g N_1_X158/M6_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX158/M8 N_X158/14_X158/M8_d N_5_X158/M8_g X158/18 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX158/M9 N_1_X158/M9_d N_35_X158/M9_g N_X158/14_X158/M8_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06 PS=1.38e-06
mX158/M10 N_X158/15_X158/M10_d N_1_X158/M10_g N_1_X158/M9_d N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06 PS=1.04e-06
mX158/M11 X158/19 N_5_X158/M11_g N_X158/15_X158/M10_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX158/M12 N_1_X158/M12_d N_X158/16_X158/M12_g X158/19 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX158/M13 X158/20 N_6_X158/M13_g N_1_X158/M12_d N_1_X154/M0_b NMOS_VTL L=5e-08
+ W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX158/M14 N_X158/16_X158/M14_d N_1_X158/M14_g X158/20 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX158/M15 N_1_X158/M15_d N_X158/16_X158/M15_g N_1_X158/M15_s N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX158/M16 N_5_X158/M16_d N_X158/CLK_X158/M16_g N_1_X158/M16_s N_5_X158/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX158/M17 N_X158/11_X158/M17_d N_X158/D_X158/M17_g N_5_X158/M16_d N_5_X158/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX158/M18 N_X158/13_X158/M18_d N_35_X158/M18_g N_X158/11_X158/M17_d
+ N_5_X158/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14 PD=1.09e-06
+ PS=1.28e-06
mX158/M19 N_X158/12_X158/M19_d N_1_X158/M19_g N_X158/13_X158/M18_d
+ N_5_X158/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14 PD=1.38e-06
+ PS=1.09e-06
mX158/M20 N_5_X158/M20_d N_1_X158/M20_g N_35_X158/M20_s N_5_X158/M16_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX158/M21 N_5_X158/M21_d N_6_X158/M21_g N_X158/12_X158/M19_d N_5_X158/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX158/M22 N_X158/12_X158/M22_d N_X158/14_X158/M22_g N_5_X158/M21_d
+ N_5_X158/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13 PD=1.21e-06
+ PS=2.33e-06
mX158/M23 N_X158/14_X158/M23_d N_5_X158/M23_g N_5_X158/M23_s N_5_X158/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX158/M24 N_1_X158/M24_d N_1_X158/M24_g N_X158/14_X158/M23_d N_5_X158/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13 PD=7.8e-07 PS=3.12e-06
mX158/M25 N_5_X158/M25_d N_X158/13_X158/M25_g N_X158/14_X158/M23_d
+ N_5_X158/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX158/M26 N_X158/15_X158/M26_d N_35_X158/M26_g N_1_X158/M24_d N_5_X158/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14 PD=3.3e-06 PS=7.8e-07
mX158/M27 N_X158/15_X158/M26_d N_X158/16_X158/M27_g N_5_X158/M25_d
+ N_5_X158/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX158/M28 N_5_X158/M28_d N_5_X158/M28_g N_X158/15_X158/M26_d N_5_X158/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX158/M29 N_X158/16_X158/M29_d N_6_X158/M29_g N_5_X158/M28_d N_5_X158/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX158/M30 N_5_X158/M30_d N_1_X158/M30_g N_X158/16_X158/M29_d N_5_X158/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06 PS=1.28e-06
mX158/M31 N_1_X158/M31_d N_X158/16_X158/M31_g N_5_X158/M30_d N_5_X158/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
mX159/M0 N_1_X159/M0_s N_X159/CLK_X159/M0_g N_1_X159/M0_s N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX159/M1 N_X159/11_X159/M1_d N_X159/D_X159/M1_g N_1_X159/M0_s N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX159/M2 N_5_X159/M2_d N_1_X159/M2_g N_1_X159/M2_s N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX159/M3 N_X159/13_X159/M3_d N_1_X159/M3_g N_X159/11_X159/M1_d N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06 PS=9.2e-07
mX159/M4 N_X159/12_X159/M4_d N_5_X159/M4_g N_X159/13_X159/M3_d N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06 PS=1.2e-06
mX159/M5 X159/17 N_6_X159/M5_g N_X159/12_X159/M4_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX159/M6 N_1_X159/M6_d N_X159/14_X159/M6_g X159/17 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX159/M7 X159/18 N_X159/13_X159/M7_g N_1_X159/M6_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX159/M8 N_X159/14_X159/M8_d N_5_X159/M8_g X159/18 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX159/M9 N_36_X159/M9_d N_5_X159/M9_g N_X159/14_X159/M8_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06 PS=1.38e-06
mX159/M10 N_X159/15_X159/M10_d N_1_X159/M10_g N_36_X159/M9_d N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06 PS=1.04e-06
mX159/M11 X159/19 N_5_X159/M11_g N_X159/15_X159/M10_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX159/M12 N_1_X159/M12_d N_X159/16_X159/M12_g X159/19 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX159/M13 X159/20 N_6_X159/M13_g N_1_X159/M12_d N_1_X154/M0_b NMOS_VTL L=5e-08
+ W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX159/M14 N_X159/16_X159/M14_d N_36_X159/M14_g X159/20 N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX159/M15 N_37_X159/M15_d N_X159/16_X159/M15_g N_1_X159/M15_s N_1_X154/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX159/M16 N_5_X159/M16_d N_X159/CLK_X159/M16_g N_1_X159/M16_s N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX159/M17 N_X159/11_X159/M17_d N_X159/D_X159/M17_g N_5_X159/M16_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX159/M18 N_X159/13_X159/M18_d N_5_X159/M18_g N_X159/11_X159/M17_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14 PD=1.09e-06
+ PS=1.28e-06
mX159/M19 N_X159/12_X159/M19_d N_1_X159/M19_g N_X159/13_X159/M18_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14 PD=1.38e-06
+ PS=1.09e-06
mX159/M20 N_5_X159/M20_d N_1_X159/M20_g N_5_X159/M20_s N_5_X153/M16_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX159/M21 N_5_X159/M21_d N_6_X159/M21_g N_X159/12_X159/M19_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX159/M22 N_X159/12_X159/M22_d N_X159/14_X159/M22_g N_5_X159/M21_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13 PD=1.21e-06
+ PS=2.33e-06
mX159/M23 N_X159/14_X159/M23_d N_5_X159/M23_g N_5_X159/M23_s N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX159/M24 N_36_X159/M24_d N_1_X159/M24_g N_X159/14_X159/M23_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13 PD=7.8e-07 PS=3.12e-06
mX159/M25 N_5_X159/M25_d N_X159/13_X159/M25_g N_X159/14_X159/M23_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX159/M26 N_X159/15_X159/M26_d N_5_X159/M26_g N_36_X159/M24_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14 PD=3.3e-06 PS=7.8e-07
mX159/M27 N_X159/15_X159/M26_d N_X159/16_X159/M27_g N_5_X159/M25_d
+ N_5_X153/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX159/M28 N_5_X159/M28_d N_5_X159/M28_g N_X159/15_X159/M26_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX159/M29 N_X159/16_X159/M29_d N_6_X159/M29_g N_5_X159/M28_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX159/M30 N_5_X159/M30_d N_36_X159/M30_g N_X159/16_X159/M29_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06 PS=1.28e-06
mX159/M31 N_37_X159/M31_d N_X159/16_X159/M31_g N_5_X159/M30_d N_5_X153/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
mX160/M0 N_1_X160/M0_s N_X160/CLK_X160/M0_g N_1_X160/M0_s N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=5.25e-14 AS=2.625e-14 PD=9.2e-07 PS=7.1e-07
mX160/M1 N_X160/11_X160/M1_d N_X160/D_X160/M1_g N_1_X160/M0_s N_1_X156/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=5.25e-14 PD=9.2e-07 PS=9.2e-07
mX160/M2 N_38_X160/M2_d N_1_X160/M2_g N_1_X160/M2_s N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.5e-14 PD=7.1e-07 PS=8.6e-07
mX160/M3 N_X160/13_X160/M3_d N_1_X160/M3_g N_X160/11_X160/M1_d N_1_X156/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=8.75e-14 AS=5.25e-14 PD=1.2e-06 PS=9.2e-07
mX160/M4 N_X160/12_X160/M4_d N_38_X160/M4_g N_X160/13_X160/M3_d N_1_X156/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=8.75e-14 PD=1.28e-06 PS=1.2e-06
mX160/M5 X160/17 N_14_X160/M5_g N_X160/12_X160/M4_d N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX160/M6 N_1_X160/M6_d N_X160/14_X160/M6_g X160/17 N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=1.8e-13 AS=7e-14 PD=1.72e-06 PS=1.28e-06
mX160/M7 X160/18 N_X160/13_X160/M7_g N_1_X160/M6_d N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=1.8e-13 PD=1.28e-06 PS=1.72e-06
mX160/M8 N_X160/14_X160/M8_d N_5_X160/M8_g X160/18 N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7.375e-14 AS=7e-14 PD=1.38e-06 PS=1.28e-06
mX160/M9 N_1_X160/M9_d N_38_X160/M9_g N_X160/14_X160/M8_d N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=6.75e-14 AS=7.375e-14 PD=1.04e-06 PS=1.38e-06
mX160/M10 N_X160/15_X160/M10_d N_1_X160/M10_g N_1_X160/M9_d N_1_X156/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=5.25e-14 AS=6.75e-14 PD=1.28e-06 PS=1.04e-06
mX160/M11 X160/19 N_5_X160/M11_g N_X160/15_X160/M10_d N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=5.25e-14 PD=1.28e-06 PS=1.28e-06
mX160/M12 N_1_X160/M12_d N_X160/16_X160/M12_g X160/19 N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=9e-14 AS=7e-14 PD=1.36e-06 PS=1.28e-06
mX160/M13 X160/20 N_14_X160/M13_g N_1_X160/M12_d N_1_X156/M0_b NMOS_VTL L=5e-08
+ W=5e-07 AD=7e-14 AS=9e-14 PD=1.28e-06 PS=1.36e-06
mX160/M14 N_X160/16_X160/M14_d N_1_X160/M14_g X160/20 N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=4.64625e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX160/M15 N_1_X160/M15_d N_X160/16_X160/M15_g N_1_X160/M15_s N_1_X156/M0_b
+ NMOS_VTL L=5e-08 W=2.5e-07 AD=2.625e-14 AS=4.115e-14 PD=7.1e-07 PS=8.6e-07
mX160/M16 N_5_X160/M16_d N_X160/CLK_X160/M16_g N_1_X160/M16_s N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.075e-13 AS=5.25e-14 PD=1.43e-06 PS=1.21e-06
mX160/M17 N_X160/11_X160/M17_d N_X160/D_X160/M17_g N_5_X160/M16_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.075e-13 PD=1.28e-06 PS=1.43e-06
mX160/M18 N_X160/13_X160/M18_d N_38_X160/M18_g N_X160/11_X160/M17_d
+ N_5_X156/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=7.375e-14 AS=5.25e-14 PD=1.09e-06
+ PS=1.28e-06
mX160/M19 N_X160/12_X160/M19_d N_1_X160/M19_g N_X160/13_X160/M18_d
+ N_5_X156/M16_b PMOS_VTL L=5e-08 W=2.5e-07 AD=6.5e-14 AS=7.375e-14 PD=1.38e-06
+ PS=1.09e-06
mX160/M20 N_5_X160/M20_d N_1_X160/M20_g N_38_X160/M20_s N_5_X156/M16_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX160/M21 N_5_X160/M21_d N_14_X160/M21_g N_X160/12_X160/M19_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.5415e-13 AS=6.5e-14 PD=2.33e-06 PS=1.38e-06
mX160/M22 N_X160/12_X160/M22_d N_X160/14_X160/M22_g N_5_X160/M21_d
+ N_5_X156/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.5415e-13 PD=1.21e-06
+ PS=2.33e-06
mX160/M23 N_X160/14_X160/M23_d N_5_X160/M23_g N_5_X160/M23_s N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.9415e-13 AS=9.7675e-14 PD=3.12e-06 PS=1.895e-06
mX160/M24 N_1_X160/M24_d N_1_X160/M24_g N_X160/14_X160/M23_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.5e-14 AS=1.9415e-13 PD=7.8e-07 PS=3.12e-06
mX160/M25 N_5_X160/M25_d N_X160/13_X160/M25_g N_X160/14_X160/M23_d
+ N_5_X156/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.9415e-13 PD=1.28e-06
+ PS=3.12e-06
mX160/M26 N_X160/15_X160/M26_d N_38_X160/M26_g N_1_X160/M24_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=2.5e-07 AD=3.058e-13 AS=3.5e-14 PD=3.3e-06 PS=7.8e-07
mX160/M27 N_X160/15_X160/M26_d N_X160/16_X160/M27_g N_5_X160/M25_d
+ N_5_X156/M16_b PMOS_VTL L=5e-08 W=5e-07 AD=3.058e-13 AS=7e-14 PD=3.3e-06
+ PS=1.28e-06
mX160/M28 N_5_X160/M28_d N_5_X160/M28_g N_X160/15_X160/M26_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.22675e-13 AS=3.058e-13 PD=1.995e-06 PS=3.3e-06
mX160/M29 N_X160/16_X160/M29_d N_14_X160/M29_g N_5_X160/M28_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=7e-14 AS=1.22675e-13 PD=1.28e-06 PS=1.995e-06
mX160/M30 N_5_X160/M30_d N_1_X160/M30_g N_X160/16_X160/M29_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=1.025e-13 AS=7e-14 PD=1.41e-06 PS=1.28e-06
mX160/M31 N_1_X160/M31_d N_X160/16_X160/M31_g N_5_X160/M30_d N_5_X156/M16_b
+ PMOS_VTL L=5e-08 W=5e-07 AD=5.25e-14 AS=1.025e-13 PD=1.21e-06 PS=1.41e-06
mX161/M0 N_12_X161/M0_d N_12_X161/M0_g N_1_X161/M0_s N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=6.675e-07 AD=9.345e-14 AS=2.2695e-13 PD=1.615e-06 PS=2.015e-06
mX161/M1 N_1_X161/M1_d N_12_X161/M1_g N_12_X161/M0_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=6.675e-07 AD=9.3275e-14 AS=9.345e-14 PD=1.615e-06 PS=1.615e-06
mX161/M2 N_12_X161/M2_d N_12_X161/M2_g N_1_X161/M1_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=6.65e-07 AD=6.9825e-14 AS=9.3275e-14 PD=1.54e-06 PS=1.615e-06
mX161/M3 N_12_X161/M3_d N_12_X161/M3_g N_5_X161/M3_s N_5_X158/M16_b PMOS_VTL
+ L=5e-08 W=1e-06 AD=1.4e-13 AS=3.4e-13 PD=2.28e-06 PS=2.68e-06
mX161/M4 N_5_X161/M4_d N_12_X161/M4_g N_12_X161/M3_d N_5_X158/M16_b PMOS_VTL
+ L=5e-08 W=1e-06 AD=1.4e-13 AS=1.4e-13 PD=2.28e-06 PS=2.28e-06
mX161/M5 N_12_X161/M5_d N_12_X161/M5_g N_5_X161/M4_d N_5_X158/M16_b PMOS_VTL
+ L=5e-08 W=1e-06 AD=1.4e-13 AS=1.4e-13 PD=2.28e-06 PS=2.28e-06
mX161/M6 N_5_X161/M6_d N_12_X161/M6_g N_12_X161/M5_d N_5_X158/M16_b PMOS_VTL
+ L=5e-08 W=1e-06 AD=1.05e-13 AS=1.4e-13 PD=2.21e-06 PS=2.28e-06
mX162/M0 N_39_X162/M0_d N_15_X162/M0_g N_1_X162/M0_s N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=6.675e-07 AD=9.345e-14 AS=2.2695e-13 PD=1.615e-06 PS=2.015e-06
mX162/M1 N_1_X162/M1_d N_15_X162/M1_g N_39_X162/M0_d N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=6.675e-07 AD=9.3275e-14 AS=9.345e-14 PD=1.615e-06 PS=1.615e-06
mX162/M2 N_39_X162/M2_d N_15_X162/M2_g N_1_X162/M1_d N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=6.65e-07 AD=6.9825e-14 AS=9.3275e-14 PD=1.54e-06 PS=1.615e-06
mX162/M3 N_39_X162/M3_d N_15_X162/M3_g N_5_X162/M3_s N_5_X162/M3_b PMOS_VTL
+ L=5e-08 W=1e-06 AD=1.4e-13 AS=3.4e-13 PD=2.28e-06 PS=2.68e-06
mX162/M4 N_5_X162/M4_d N_15_X162/M4_g N_39_X162/M3_d N_5_X162/M3_b PMOS_VTL
+ L=5e-08 W=1e-06 AD=1.4e-13 AS=1.4e-13 PD=2.28e-06 PS=2.28e-06
mX162/M5 N_39_X162/M5_d N_15_X162/M5_g N_5_X162/M4_d N_5_X162/M3_b PMOS_VTL
+ L=5e-08 W=1e-06 AD=1.4e-13 AS=1.4e-13 PD=2.28e-06 PS=2.28e-06
mX162/M6 N_5_X162/M6_d N_15_X162/M6_g N_39_X162/M5_d N_5_X162/M3_b PMOS_VTL
+ L=5e-08 W=1e-06 AD=1.05e-13 AS=1.4e-13 PD=2.21e-06 PS=2.28e-06
mX163/M0 N_1_X163/M0_d N_X163/A_X163/M0_g N_1_X163/M0_s N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX163/M1 N_1_X163/M1_d N_X163/A_X163/M1_g N_5_X163/M1_s N_5_X158/M16_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX164/M0 N_9_X164/M0_d N_X164/A_X164/M0_g N_1_X164/M0_s N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX164/M1 N_9_X164/M1_d N_X164/A_X164/M1_g N_5_X164/M1_s N_5_X156/M16_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX165/M0 N_8_X165/M0_d N_X165/A_X165/M0_g N_1_X165/M0_s N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX165/M1 N_8_X165/M1_d N_X165/A_X165/M1_g N_5_X165/M1_s N_5_X162/M3_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX166/M0 N_14_X166/M0_d N_X166/A_X166/M0_g N_1_X166/M0_s N_1_X156/M0_b NMOS_VTL
+ L=5e-08 W=2.5e-07 AD=2.625e-14 AS=2.625e-14 PD=7.1e-07 PS=7.1e-07
mX166/M1 N_14_X166/M1_d N_X166/A_X166/M1_g N_5_X166/M1_s N_5_X162/M3_b PMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=5.25e-14 PD=1.21e-06 PS=1.21e-06
mX167/M0 N_1_X167/M0_d N_40_X167/M0_g N_1_X167/M0_s N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=8.75e-14 PD=1.28e-06 PS=1.35e-06
mX167/M1 N_1_X167/M1_d N_40_X167/M1_g N_1_X167/M0_d N_1_X154/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX167/M2 N_1_X167/M2_d N_40_X167/M2_g N_5_X167/M2_s N_5_X153/M16_b PMOS_VTL
+ L=5e-08 W=1e-06 AD=1.4e-13 AS=1.05e-13 PD=2.28e-06 PS=2.21e-06
mX167/M3 N_5_X167/M3_d N_40_X167/M3_g N_1_X167/M2_d N_5_X153/M16_b PMOS_VTL
+ L=5e-08 W=1e-06 AD=1.05e-13 AS=1.4e-13 PD=2.21e-06 PS=2.28e-06
mX168/M0 N_41_X168/M0_d N_1_X168/M0_g N_1_X168/M0_s N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=7e-14 AS=8.75e-14 PD=1.28e-06 PS=1.35e-06
mX168/M1 N_1_X168/M1_d N_1_X168/M1_g N_41_X168/M0_d N_1_X153/M0_b NMOS_VTL
+ L=5e-08 W=5e-07 AD=5.25e-14 AS=7e-14 PD=1.21e-06 PS=1.28e-06
mX168/M2 N_41_X168/M2_d N_1_X168/M2_g N_5_X168/M2_s N_5_X156/M16_b PMOS_VTL
+ L=5e-08 W=1e-06 AD=1.4e-13 AS=1.05e-13 PD=2.28e-06 PS=2.21e-06
mX168/M3 N_5_X168/M3_d N_1_X168/M3_g N_41_X168/M2_d N_5_X156/M16_b PMOS_VTL
+ L=5e-08 W=1e-06 AD=1.05e-13 AS=1.4e-13 PD=2.21e-06 PS=2.28e-06
*
.include "/media/ntfsdrive1/workspace/ProjectDIC2/runsets/pex/extracted.sp.FULLSYSTEM.pxi"
*
.ends
*
*
