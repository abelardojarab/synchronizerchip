module XOR2X1 (
	Y, 
	B, 
	A);
   output Y;
   input B;
   input A;
endmodule

module OR2X1 (
	Y, 
	B, 
	A);
   output Y;
   input B;
   input A;
endmodule

module NOR2X1 (
	Y, 
	B, 
	A);
   output Y;
   input B;
   input A;
endmodule

module INVX8 (
	Y, 
	A);
   output Y;
   input A;
endmodule

module INVX4 (
	Y, 
	A);
   output Y;
   input A;
endmodule

module INVX1 (
	Y, 
	A);
   output Y;
   input A;
endmodule

module FILL ();
endmodule

module DFFSR (
	S, 
	R, 
	Q, 
	D, 
	CLK);
   input S;
   input R;
   output Q;
   input D;
   input CLK;
endmodule

module BUFX2 (
	Y, 
	A);
   output Y;
   input A;
endmodule

module AOI22X1 (
	Y, 
	D, 
	C, 
	B, 
	A);
   output Y;
   input D;
   input C;
   input B;
   input A;
endmodule

module AND2X1 (
	Y, 
	B, 
	A);
   output Y;
   input B;
   input A;
endmodule

