** Generated for: hspiceD
** Generated on: Dec  9 13:43:48 2015
** Design library name: fullsystem
** Design cell name: fullsystem_tb
** Design view name: schematic
.GLOBAL vdd!


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: freepdk45_cells
** Cell name: NOR2X1
** View name: schematic
.subckt NOR2X1 a b y gnd vdd
m2 y a gnd gnd NMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
m3 gnd b y gnd NMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
m1 y b a_9_54__ vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
m0 a_9_54__ a vdd vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
.ends NOR2X1
** End of subcircuit definition.

** Library name: freepdk45_cells
** Cell name: XOR2X1
** View name: schematic
.subckt XOR2X1 a b y gnd vdd
m2 y a a_18_54__ vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
m1 a_18_54__ a_13_43__ vdd vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
m3 a_35_54__ a_2_6__ y vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
m4 vdd b a_35_54__ vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
m0 vdd a a_2_6__ vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
m5 a_13_43__ b vdd vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
m8 y a_2_6__ a_18_6__ gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m7 a_18_6__ a_13_43__ gnd gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m9 a_35_6__ a y gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m10 gnd b a_35_6__ gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m6 gnd a a_2_6__ gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m11 a_13_43__ b gnd gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
.ends XOR2X1
** End of subcircuit definition.

** Library name: fullsystem
** Cell name: DFFSR
** View name: schematic
.subckt DFFSR clk d q r s
m6 vdd d a_57_6__ vdd PMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m8 a_47_71__ clk vdd vdd PMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m15 vdd a_122_6__ q vdd PMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m0 a_2_6__ r vdd vdd PMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m1 vdd a_10_61__ a_2_6__ vdd PMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m12 vdd r a_122_6__ vdd PMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m11 a_122_6__ a_105_6__ vdd vdd PMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m4 a_23_27__ a_47_71__ a_2_6__ vdd PMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
m2 a_10_61__ a_23_27__ vdd vdd PMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m7 vdd a_47_71__ a_47_4__ vdd PMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m9 a_105_6__ a_47_71__ a_10_61__ vdd PMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
m3 vdd s a_10_61__ vdd PMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m5 a_57_6__ a_47_4__ a_23_27__ vdd PMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
m10 a_113_6__ a_47_4__ a_105_6__ vdd PMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
m13 a_113_6__ a_122_6__ vdd vdd PMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m14 vdd s a_113_6__ vdd PMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m16 a_10_6__ r a_2_6__ gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m17 gnd a_10_61__ a_10_6__ gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m28 gnd r a_130_6__ gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m27 a_130_6__ a_105_6__ a_122_6__ gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m18 a_26_6__ a_23_27__ gnd gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m19 a_10_61__ s a_26_6__ gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m30 a_113_6__ s a_146_6__ gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m29 a_146_6__ a_122_6__ gnd gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m22 gnd d a_57_6__ gnd NMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
m24 a_47_71__ clk gnd gnd NMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
m31 gnd a_122_6__ q gnd NMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
m25 a_105_6__ a_47_4__ a_10_61__ gnd NMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
m20 a_23_27__ a_47_4__ a_2_6__ gnd NMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
m23 gnd a_47_71__ a_47_4__ gnd NMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
m21 a_57_6__ a_47_71__ a_23_27__ gnd NMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
m26 a_113_6__ a_47_71__ a_105_6__ gnd NMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
.ends DFFSR
** End of subcircuit definition.

** Library name: freepdk45_cells
** Cell name: INVX1
** View name: schematic
.subckt INVX1 a y gnd vdd
m0 y a vdd vdd PMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m1 y a gnd gnd NMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
.ends INVX1
** End of subcircuit definition.

** Library name: freepdk45_cells
** Cell name: AND2X2
** View name: schematic
.subckt AND2X2 a b y gnd vdd
m0 a_2_6__ a vdd vdd PMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m1 vdd b a_2_6__ vdd PMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m2 y a_2_6__ vdd vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
m3 a_9_6__ a a_2_6__ gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m4 gnd b a_9_6__ gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m5 y a_2_6__ gnd gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
.ends AND2X2
** End of subcircuit definition.

** Library name: fullsystem
** Cell name: AOI22X1
** View name: schematic
.subckt AOI22X1 a b c d y
m5 y b a_11_6__ gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m4 a_11_6__ a gnd gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m7 gnd c a_28_6__ gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m6 a_28_6__ d y gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
m1 a_2_54__ b vdd vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
m0 vdd a a_2_54__ vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
m2 y d a_2_54__ vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
m3 a_2_54__ c y vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
.ends AOI22X1
** End of subcircuit definition.

** Library name: freepdk45_cells
** Cell name: OR2X2
** View name: schematic
.subckt OR2X2 a b y gnd vdd
m0 a_9_54__ a a_2_54__ vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
m1 vdd b a_9_54__ vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
m2 y a_2_54__ vdd vdd PMOS_VTL L=50e-9 W=1e-6 AD=0 AS=0 PD=0 PS=0 M=1
m4 gnd b a_2_54__ gnd NMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
m3 a_2_54__ a gnd gnd NMOS_VTL L=50e-9 W=250e-9 AD=0 AS=0 PD=0 PS=0 M=1
m5 y a_2_54__ gnd gnd NMOS_VTL L=50e-9 W=500e-9 AD=0 AS=0 PD=0 PS=0 M=1
.ends OR2X2
** End of subcircuit definition.

** Library name: fullsystem
** Cell name: fullsystem
** View name: schematic
.subckt fullsystem clk1 clk2 reset1 reset2 start ready rcv
xtalker_str_1xfsm_unitxu12 talker_str_1xfsm_unitxstate_regx0x talker_str_1xfsm_unitxn8 ready net70 net71 NOR2X1
xtalker_str_1xfsm_unitxu13 talker_str_1xfsm_unitxstate_regx1x talker_str_1xfsm_unitxstate_regx0x talker_str_1xfsm_unitxn8 net72 net73 XOR2X1
xtalker_str_1xsync_unitxmeta_reg_reg clk2 n19 talker_str_1xsync_unitxmeta_reg talker_str_1xfsm_unitxn4 vdd! DFFSR
xtalker_str_1xsync_unitxsync_reg_reg clk2 n16 rcv talker_str_1xfsm_unitxn4 vdd! DFFSR
xlistener_str_1xsync_unitxsync_reg_reg clk1 n22 listener_str_1xreq_sync listener_str_1xsync_unitxn2 vdd! DFFSR
xlistener_str_1xfsm_unitxack_buf_reg_reg clk1 n25 ack_out listener_str_1xsync_unitxn2 vdd! DFFSR
xlistener_str_1xsync_unitxmeta_reg_reg clk1 n28 listener_str_1xsync_unitxmeta_reg listener_str_1xsync_unitxn2 vdd! DFFSR
xtalker_str_1xfsm_unitxreq_buf_reg_reg clk2 n7 req_in talker_str_1xfsm_unitxn4 vdd! DFFSR
xtalker_str_1xfsm_unitxstate_reg_regx1x clk2 talker_str_1xfsm_unitxstate_nextx1x talker_str_1xfsm_unitxstate_regx1x talker_str_1xfsm_unitxn4 vdd! DFFSR
xtalker_str_1xfsm_unitxstate_reg_regx0x clk2 n7 talker_str_1xfsm_unitxstate_regx0x talker_str_1xfsm_unitxn4 vdd! DFFSR
xu13 rcv talker_str_1xfsm_unitxn7 net74 net75 INVX1
xu8 n6 n7 net76 net77 INVX1
xu14 talker_str_1xfsm_unitxstate_regx0x talker_str_1xfsm_unitxn6 net78 net79 INVX1
xu6 n18 n19 net80 net81 INVX1
xu5 ack_out n18 net82 net83 INVX1
xu2 talker_str_1xsync_unitxmeta_reg n15 net84 net85 INVX1
xu3 n15 n16 net86 net87 INVX1
xu20 n24 n25 net88 net89 INVX1
xu19 listener_str_1xreq_sync n24 net90 net91 INVX1
xu17 n21 n22 net92 net93 INVX1
xu23 n27 n28 net94 net95 INVX1
xu22 req_in n27 net96 net97 INVX1
xu16 listener_str_1xsync_unitxmeta_reg n21 net98 net99 INVX1
xtalker_str_1xfsm_unitxu5 reset2 talker_str_1xfsm_unitxn4 net100 net101 INVX1
xlistener_str_1xsync_unitxu4 reset1 listener_str_1xsync_unitxn2 net102 net103 INVX1
xu7 rcv talker_str_1xfsm_unitxn8 talker_str_1xfsm_unitxstate_nextx1x net104 net105 AND2X2
xtalker_str_1xfsm_unitxu11 talker_str_1xfsm_unitxstate_regx0x talker_str_1xfsm_unitxn7 start talker_str_1xfsm_unitxn6 talker_str_1xfsm_unitxn9 AOI22X1
xu1 talker_str_1xfsm_unitxstate_regx1x talker_str_1xfsm_unitxn9 n6 net106 net107 OR2X2
.ends fullsystem
** End of subcircuit definition.

** Library name: fullsystem
** Cell name: fullsystem_tb
** View name: schematic
xfullsystem net7 net6 net5 net4 net3 net2 net1 fullsystem
.END
